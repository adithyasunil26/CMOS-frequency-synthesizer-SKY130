magic
tech sky130A
magscale 1 2
timestamp 1640805170
<< ndiff >>
rect 1840 -30 1980 110
rect 2720 92 2860 110
rect 2720 -8 2740 92
rect 2840 -8 2860 92
rect 2720 -30 2860 -8
rect 3600 92 3740 110
rect 3600 -8 3620 92
rect 3720 -8 3740 92
rect 3600 -30 3740 -8
rect 4460 92 4600 110
rect 4460 -8 4480 92
rect 4580 -8 4600 92
rect 4460 -30 4600 -8
rect 5320 92 5460 110
rect 5320 -8 5340 92
rect 5440 -8 5460 92
rect 5320 -30 5460 -8
rect 6220 92 6360 110
rect 6220 -8 6240 92
rect 6340 -8 6360 92
rect 6220 -30 6360 -8
<< ndiffc >>
rect 2740 -8 2840 92
rect 3620 -8 3720 92
rect 4480 -8 4580 92
rect 5340 -8 5440 92
rect 6240 -8 6340 92
<< psubdiff >>
rect 4650 -1430 4910 -1400
rect 4650 -1630 4680 -1430
rect 4880 -1630 4910 -1430
rect 4650 -1660 4910 -1630
<< psubdiffcont >>
rect 4680 -1630 4880 -1430
<< locali >>
rect 300 1520 490 1540
rect 300 1390 320 1520
rect 270 1370 320 1390
rect 470 1370 490 1520
rect 270 1350 490 1370
rect 2110 190 2120 260
rect 2990 190 3000 260
rect 3870 190 3880 260
rect 4730 190 4740 260
rect 5590 190 5600 260
rect 6490 190 6500 260
rect 1840 90 1980 110
rect 1840 -10 1860 90
rect 1960 -10 1980 90
rect 1840 -30 1980 -10
rect 2720 92 2860 110
rect 2720 -10 2740 92
rect 2840 -10 2860 92
rect 2720 -30 2860 -10
rect 3600 92 3740 110
rect 3600 -10 3620 92
rect 3720 -10 3740 92
rect 3600 -30 3740 -10
rect 4460 92 4600 110
rect 4460 -10 4480 92
rect 4580 -10 4600 92
rect 4460 -30 4600 -10
rect 5320 92 5460 110
rect 5320 -10 5340 92
rect 5440 -10 5460 92
rect 5320 -30 5460 -10
rect 6220 92 6360 110
rect 6220 -10 6240 92
rect 6340 -10 6360 92
rect 6220 -30 6360 -10
rect 730 -190 970 -170
rect 730 -390 750 -190
rect 950 -390 970 -190
rect 730 -410 970 -390
rect 2110 -1410 2210 -1270
rect 2990 -1410 3090 -1280
rect 3870 -1410 3970 -1280
rect 4730 -1410 4830 -1280
rect 5590 -1410 5690 -1280
rect 6490 -1410 6590 -1280
rect 2040 -1430 2280 -1410
rect 2040 -1630 2060 -1430
rect 2260 -1630 2280 -1430
rect 2040 -1650 2280 -1630
rect 2920 -1430 3160 -1410
rect 2920 -1630 2940 -1430
rect 3140 -1630 3160 -1430
rect 2920 -1650 3160 -1630
rect 3800 -1430 4040 -1410
rect 3800 -1630 3820 -1430
rect 4020 -1630 4040 -1430
rect 3800 -1650 4040 -1630
rect 4660 -1430 4900 -1410
rect 4660 -1630 4680 -1430
rect 4880 -1630 4900 -1430
rect 4660 -1650 4900 -1630
rect 5520 -1430 5760 -1410
rect 5520 -1630 5540 -1430
rect 5740 -1630 5760 -1430
rect 5520 -1650 5760 -1630
rect 6430 -1430 6670 -1410
rect 6430 -1630 6450 -1430
rect 6650 -1630 6670 -1430
rect 6430 -1650 6670 -1630
<< viali >>
rect 320 1370 470 1520
rect 1860 -10 1960 90
rect 2740 -8 2840 90
rect 2740 -10 2840 -8
rect 3620 -8 3720 90
rect 3620 -10 3720 -8
rect 4480 -8 4580 90
rect 4480 -10 4580 -8
rect 5340 -8 5440 90
rect 5340 -10 5440 -8
rect 6240 -8 6340 90
rect 6240 -10 6340 -8
rect 750 -390 950 -190
rect 2060 -1630 2260 -1430
rect 2940 -1630 3140 -1430
rect 3820 -1630 4020 -1430
rect 4680 -1630 4880 -1430
rect 5540 -1630 5740 -1430
rect 6450 -1630 6650 -1430
<< metal1 >>
rect 300 1520 490 1540
rect 300 1370 320 1520
rect 470 1370 490 1520
rect 300 1350 490 1370
rect 1840 90 1980 110
rect 1840 -10 1860 90
rect 1960 -10 1980 90
rect 1840 -30 1980 -10
rect 2720 90 2860 110
rect 2720 -10 2740 90
rect 2840 -10 2860 90
rect 2720 -30 2860 -10
rect 3600 90 3740 110
rect 3600 -10 3620 90
rect 3720 -10 3740 90
rect 3600 -30 3740 -10
rect 4460 90 4600 110
rect 4460 -10 4480 90
rect 4580 -10 4600 90
rect 4460 -30 4600 -10
rect 5320 90 5460 110
rect 5320 -10 5340 90
rect 5440 -10 5460 90
rect 5320 -30 5460 -10
rect 6220 90 6360 110
rect 6220 -10 6240 90
rect 6340 -10 6360 90
rect 6220 -30 6360 -10
rect 730 -190 970 -170
rect 730 -390 750 -190
rect 950 -390 970 -190
rect 730 -410 970 -390
rect 2040 -1430 2280 -1410
rect 2040 -1630 2060 -1430
rect 2260 -1630 2280 -1430
rect 2040 -1650 2280 -1630
rect 2920 -1430 3160 -1410
rect 2920 -1630 2940 -1430
rect 3140 -1630 3160 -1430
rect 2920 -1650 3160 -1630
rect 3800 -1430 4040 -1410
rect 3800 -1630 3820 -1430
rect 4020 -1630 4040 -1430
rect 3800 -1650 4040 -1630
rect 4660 -1430 4900 -1410
rect 4660 -1630 4680 -1430
rect 4880 -1630 4900 -1430
rect 4660 -1650 4900 -1630
rect 5520 -1430 5760 -1410
rect 5520 -1630 5540 -1430
rect 5740 -1630 5760 -1430
rect 5520 -1650 5760 -1630
rect 6430 -1430 6670 -1410
rect 6430 -1630 6450 -1430
rect 6650 -1630 6670 -1430
rect 6430 -1650 6670 -1630
<< via1 >>
rect 320 1370 470 1520
rect 1860 -10 1960 90
rect 2740 -10 2840 90
rect 3620 -10 3720 90
rect 4480 -10 4580 90
rect 5340 -10 5440 90
rect 6240 -10 6340 90
rect 750 -390 950 -190
rect 2060 -1630 2260 -1430
rect 2940 -1630 3140 -1430
rect 3820 -1630 4020 -1430
rect 4680 -1630 4880 -1430
rect 5540 -1630 5740 -1430
rect 6450 -1630 6650 -1430
<< metal2 >>
rect 300 1520 490 1540
rect 300 1370 320 1520
rect 470 1370 490 1520
rect 300 1350 490 1370
rect 1840 90 1980 110
rect 1840 -10 1860 90
rect 1960 -10 1980 90
rect 1840 -30 1980 -10
rect 2720 90 2860 110
rect 2720 -10 2740 90
rect 2840 -10 2860 90
rect 2720 -30 2860 -10
rect 3600 90 3740 110
rect 3600 -10 3620 90
rect 3720 -10 3740 90
rect 3600 -30 3740 -10
rect 4460 90 4600 110
rect 4460 -10 4480 90
rect 4580 -10 4600 90
rect 4460 -30 4600 -10
rect 5320 90 5460 110
rect 5320 -10 5340 90
rect 5440 -10 5460 90
rect 5320 -30 5460 -10
rect 6220 90 6360 110
rect 6220 -10 6240 90
rect 6340 -10 6360 90
rect 6220 -30 6360 -10
rect 730 -190 970 -170
rect 730 -390 750 -190
rect 950 -390 970 -190
rect 730 -410 970 -390
rect 2040 -1430 2280 -1410
rect 2040 -1630 2060 -1430
rect 2260 -1630 2280 -1430
rect 2040 -1650 2280 -1630
rect 2920 -1430 3160 -1410
rect 2920 -1630 2940 -1430
rect 3140 -1630 3160 -1430
rect 2920 -1650 3160 -1630
rect 3800 -1430 4040 -1410
rect 3800 -1630 3820 -1430
rect 4020 -1630 4040 -1430
rect 3800 -1650 4040 -1630
rect 4660 -1430 4900 -1410
rect 4660 -1630 4680 -1430
rect 4880 -1630 4900 -1430
rect 4660 -1650 4900 -1630
rect 5520 -1430 5760 -1410
rect 5520 -1630 5540 -1430
rect 5740 -1630 5760 -1430
rect 5520 -1650 5760 -1630
rect 6430 -1430 6670 -1410
rect 6430 -1630 6450 -1430
rect 6650 -1630 6670 -1430
rect 6430 -1650 6670 -1630
<< via2 >>
rect 320 1370 470 1520
rect 1860 -10 1960 90
rect 2740 -10 2840 90
rect 3620 -10 3720 90
rect 4480 -10 4580 90
rect 5340 -10 5440 90
rect 6240 -10 6340 90
rect 750 -390 950 -190
rect 2060 -1630 2260 -1430
rect 2940 -1630 3140 -1430
rect 3820 -1630 4020 -1430
rect 4680 -1630 4880 -1430
rect 5540 -1630 5740 -1430
rect 6450 -1630 6650 -1430
<< metal3 >>
rect 300 1520 490 1540
rect 300 1370 320 1520
rect 470 1370 490 1520
rect 300 1350 490 1370
rect 230 30 1460 1230
rect 1570 490 2320 1250
rect 2430 490 3180 1250
rect 3350 490 4100 1250
rect 4220 490 4970 1250
rect 5090 490 5840 1250
rect 5970 490 6720 1250
rect 1840 90 1980 490
rect 750 -170 950 30
rect 1840 -10 1860 90
rect 1960 -10 1980 90
rect 1840 -30 1980 -10
rect 2720 90 2860 490
rect 2720 -10 2740 90
rect 2840 -10 2860 90
rect 2720 -30 2860 -10
rect 3600 90 3740 490
rect 3600 -10 3620 90
rect 3720 -10 3740 90
rect 3600 -30 3740 -10
rect 4460 90 4600 490
rect 4460 -10 4480 90
rect 4580 -10 4600 90
rect 4460 -30 4600 -10
rect 5320 90 5460 490
rect 5320 -10 5340 90
rect 5440 -10 5460 90
rect 5320 -30 5460 -10
rect 6220 90 6360 490
rect 6220 -10 6240 90
rect 6340 -10 6360 90
rect 6220 -30 6360 -10
rect 730 -190 970 -170
rect 730 -390 750 -190
rect 950 -390 970 -190
rect 730 -410 970 -390
rect 2040 -1430 2280 -1410
rect 2040 -1630 2060 -1430
rect 2260 -1630 2280 -1430
rect 2040 -1650 2280 -1630
rect 2920 -1430 3160 -1410
rect 2920 -1630 2940 -1430
rect 3140 -1630 3160 -1430
rect 2920 -1650 3160 -1630
rect 3800 -1430 4040 -1410
rect 3800 -1630 3820 -1430
rect 4020 -1630 4040 -1430
rect 3800 -1650 4040 -1630
rect 4660 -1430 4900 -1410
rect 4660 -1630 4680 -1430
rect 4880 -1630 4900 -1430
rect 4660 -1650 4900 -1630
rect 5520 -1430 5760 -1410
rect 5520 -1630 5540 -1430
rect 5740 -1630 5760 -1430
rect 5520 -1650 5760 -1630
rect 6430 -1430 6670 -1410
rect 6430 -1630 6450 -1430
rect 6650 -1630 6670 -1430
rect 6430 -1650 6670 -1630
<< via3 >>
rect 320 1370 470 1520
rect 750 -390 950 -190
rect 2060 -1630 2260 -1430
rect 2940 -1630 3140 -1430
rect 3820 -1630 4020 -1430
rect 4680 -1630 4880 -1430
rect 5540 -1630 5740 -1430
rect 6450 -1630 6650 -1430
<< mimcap >>
rect 330 1090 1370 1130
rect 330 170 370 1090
rect 1330 170 1370 1090
rect 1670 1110 2230 1150
rect 1670 630 1710 1110
rect 2190 630 2230 1110
rect 1670 590 2230 630
rect 2530 1110 3090 1150
rect 2530 630 2570 1110
rect 3050 630 3090 1110
rect 2530 590 3090 630
rect 3450 1110 4010 1150
rect 3450 630 3490 1110
rect 3970 630 4010 1110
rect 3450 590 4010 630
rect 4320 1110 4880 1150
rect 4320 630 4360 1110
rect 4840 630 4880 1110
rect 4320 590 4880 630
rect 5190 1110 5750 1150
rect 5190 630 5230 1110
rect 5710 630 5750 1110
rect 5190 590 5750 630
rect 6070 1110 6630 1150
rect 6070 630 6110 1110
rect 6590 630 6630 1110
rect 6070 590 6630 630
rect 330 130 1370 170
<< mimcapcontact >>
rect 370 170 1330 1090
rect 1710 630 2190 1110
rect 2570 630 3050 1110
rect 3490 630 3970 1110
rect 4360 630 4840 1110
rect 5230 630 5710 1110
rect 6110 630 6590 1110
<< metal4 >>
rect 290 1520 6780 1550
rect 290 1370 320 1520
rect 470 1370 6780 1520
rect 290 1340 6780 1370
rect 630 1091 840 1340
rect 1810 1111 2010 1340
rect 2670 1111 2870 1340
rect 3590 1111 3790 1340
rect 4460 1111 4660 1340
rect 5330 1111 5530 1340
rect 6210 1111 6410 1340
rect 1709 1110 2191 1111
rect 369 1090 1331 1091
rect 369 170 370 1090
rect 1330 170 1331 1090
rect 1709 630 1710 1110
rect 2190 630 2191 1110
rect 1709 629 2191 630
rect 2569 1110 3051 1111
rect 2569 630 2570 1110
rect 3050 630 3051 1110
rect 2569 629 3051 630
rect 3489 1110 3971 1111
rect 3489 630 3490 1110
rect 3970 630 3971 1110
rect 3489 629 3971 630
rect 4359 1110 4841 1111
rect 4359 630 4360 1110
rect 4840 630 4841 1110
rect 4359 629 4841 630
rect 5229 1110 5711 1111
rect 5229 630 5230 1110
rect 5710 630 5711 1110
rect 5229 629 5711 630
rect 6109 1110 6591 1111
rect 6109 630 6110 1110
rect 6590 630 6591 1110
rect 6109 629 6591 630
rect 369 169 1331 170
rect 230 -190 1490 -140
rect 230 -390 750 -190
rect 950 -390 1490 -190
rect 230 -440 1490 -390
rect 1190 -1380 1490 -440
rect 1190 -1430 7710 -1380
rect 1190 -1630 2060 -1430
rect 2260 -1630 2940 -1430
rect 3140 -1630 3820 -1430
rect 4020 -1630 4680 -1430
rect 4880 -1630 5540 -1430
rect 5740 -1630 6450 -1430
rect 6650 -1630 7710 -1430
rect 1190 -1680 7710 -1630
use switch  switch_1
timestamp 1640608635
transform 1 0 2890 0 1 -1308
box -190 -40 240 1600
use switch  switch_0
timestamp 1640608635
transform 1 0 2010 0 1 -1308
box -190 -40 240 1600
use switch  switch_2
timestamp 1640608635
transform 1 0 3770 0 1 -1308
box -190 -40 240 1600
use switch  switch_3
timestamp 1640608635
transform 1 0 4630 0 1 -1308
box -190 -40 240 1600
use switch  switch_4
timestamp 1640608635
transform 1 0 5490 0 1 -1308
box -190 -40 240 1600
use switch  switch_5
timestamp 1640608635
transform 1 0 6390 0 1 -1308
box -190 -40 240 1600
<< labels >>
rlabel locali 4750 -1370 4751 -1370 1 gnd!
rlabel locali 280 1360 280 1360 1 v
rlabel locali 2120 220 2120 220 1 a0
rlabel locali 3000 220 3000 220 1 a1
rlabel locali 3880 210 3880 210 1 a2
rlabel locali 4740 210 4740 210 1 a3
rlabel locali 5600 200 5600 200 1 a4
rlabel locali 6500 200 6500 200 1 a5
<< end >>
