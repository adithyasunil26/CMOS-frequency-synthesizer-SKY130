magic
tech sky130A
magscale 1 2
timestamp 1640921877
<< psubdiff >>
rect -3380 530 -3120 560
rect -3380 330 -3350 530
rect -3150 330 -3120 530
rect -3380 300 -3120 330
rect -2480 530 -2220 560
rect -2480 330 -2450 530
rect -2250 330 -2220 530
rect -2480 300 -2220 330
rect -1450 530 -1190 560
rect -1450 330 -1420 530
rect -1220 330 -1190 530
rect -1450 300 -1190 330
rect -420 530 -160 560
rect -420 330 -390 530
rect -190 330 -160 530
rect -420 300 -160 330
rect 610 530 870 560
rect 610 330 640 530
rect 840 330 870 530
rect 610 300 870 330
rect 1640 530 1900 560
rect 1640 330 1670 530
rect 1870 330 1900 530
rect 1640 300 1900 330
rect 2670 530 2930 560
rect 2670 330 2700 530
rect 2900 330 2930 530
rect 2670 300 2930 330
rect 3700 530 3960 560
rect 3700 330 3730 530
rect 3930 330 3960 530
rect 3700 300 3960 330
rect 4730 530 4990 560
rect 4730 330 4760 530
rect 4960 330 4990 530
rect 4730 300 4990 330
rect 5760 530 6020 560
rect 5760 330 5790 530
rect 5990 330 6020 530
rect 5760 300 6020 330
rect 6790 530 7050 560
rect 6790 330 6820 530
rect 7020 330 7050 530
rect 6790 300 7050 330
rect 7820 530 8080 560
rect 7820 330 7850 530
rect 8050 330 8080 530
rect 7820 300 8080 330
rect 8850 530 9110 560
rect 8850 330 8880 530
rect 9080 330 9110 530
rect 8850 300 9110 330
rect 9880 530 10140 560
rect 9880 330 9910 530
rect 10110 330 10140 530
rect 9880 300 10140 330
rect 10910 530 11170 560
rect 10910 330 10940 530
rect 11140 330 11170 530
rect 10910 300 11170 330
rect 11630 530 11890 560
rect 11630 330 11660 530
rect 11860 330 11890 530
rect 11630 300 11890 330
rect 11630 -710 11890 -680
rect -3380 -740 -3120 -710
rect -3380 -940 -3350 -740
rect -3150 -940 -3120 -740
rect 11630 -910 11660 -710
rect 11860 -910 11890 -710
rect 11630 -940 11890 -910
rect -3380 -970 -3120 -940
rect 11630 -1740 11890 -1710
rect -3380 -1770 -3120 -1740
rect -3380 -1970 -3350 -1770
rect -3150 -1970 -3120 -1770
rect 11630 -1940 11660 -1740
rect 11860 -1940 11890 -1740
rect 11630 -1970 11890 -1940
rect -3380 -2000 -3120 -1970
rect -3380 -2800 -3120 -2770
rect -3380 -3000 -3350 -2800
rect -3150 -3000 -3120 -2800
rect -3380 -3030 -3120 -3000
rect -3380 -3830 -3120 -3800
rect -3380 -4030 -3350 -3830
rect -3150 -4030 -3120 -3830
rect -3380 -4060 -3120 -4030
rect -3380 -4860 -3120 -4830
rect -3380 -5060 -3350 -4860
rect -3150 -5060 -3120 -4860
rect -3380 -5090 -3120 -5060
rect 11630 -2770 11890 -2740
rect 11630 -2970 11660 -2770
rect 11860 -2970 11890 -2770
rect 11630 -3000 11890 -2970
rect 11630 -3800 11890 -3770
rect 11630 -4000 11660 -3800
rect 11860 -4000 11890 -3800
rect 11630 -4030 11890 -4000
rect 11630 -4830 11890 -4800
rect 11630 -5030 11660 -4830
rect 11860 -5030 11890 -4830
rect 11630 -5060 11890 -5030
rect 11630 -5860 11890 -5830
rect -3380 -5890 -3120 -5860
rect -3380 -6090 -3350 -5890
rect -3150 -6090 -3120 -5890
rect 11630 -6060 11660 -5860
rect 11860 -6060 11890 -5860
rect 11630 -6090 11890 -6060
rect -3380 -6120 -3120 -6090
rect 11630 -6890 11890 -6860
rect -3380 -6920 -3120 -6890
rect -3380 -7120 -3350 -6920
rect -3150 -7120 -3120 -6920
rect 11630 -7090 11660 -6890
rect 11860 -7090 11890 -6890
rect 11630 -7120 11890 -7090
rect -3380 -7150 -3120 -7120
rect 11630 -7920 11890 -7890
rect -3380 -7950 -3120 -7920
rect -3380 -8150 -3350 -7950
rect -3150 -8150 -3120 -7950
rect 11630 -8120 11660 -7920
rect 11860 -8120 11890 -7920
rect 11630 -8150 11890 -8120
rect -3380 -8180 -3120 -8150
rect 11630 -8950 11890 -8920
rect -3380 -8980 -3120 -8950
rect -3380 -9180 -3350 -8980
rect -3150 -9180 -3120 -8980
rect 11630 -9150 11660 -8950
rect 11860 -9150 11890 -8950
rect 11630 -9180 11890 -9150
rect -3380 -9210 -3120 -9180
rect 11630 -9980 11890 -9950
rect -3380 -10010 -3120 -9980
rect -3380 -10210 -3350 -10010
rect -3150 -10210 -3120 -10010
rect 11630 -10180 11660 -9980
rect 11860 -10180 11890 -9980
rect 11630 -10210 11890 -10180
rect -3380 -10240 -3120 -10210
rect 11630 -11010 11890 -10980
rect -3380 -11040 -3120 -11010
rect -3380 -11240 -3350 -11040
rect -3150 -11240 -3120 -11040
rect 11630 -11210 11660 -11010
rect 11860 -11210 11890 -11010
rect 11630 -11240 11890 -11210
rect -3380 -11270 -3120 -11240
rect 11630 -12040 11890 -12010
rect -3380 -12070 -3120 -12040
rect -3380 -12270 -3350 -12070
rect -3150 -12270 -3120 -12070
rect 11630 -12240 11660 -12040
rect 11860 -12240 11890 -12040
rect 11630 -12270 11890 -12240
rect -3380 -12300 -3120 -12270
rect 11630 -13070 11890 -13040
rect -3380 -13100 -3120 -13070
rect -3380 -13300 -3350 -13100
rect -3150 -13300 -3120 -13100
rect 11630 -13270 11660 -13070
rect 11860 -13270 11890 -13070
rect 11630 -13300 11890 -13270
rect -3380 -13330 -3120 -13300
rect 11630 -14100 11890 -14070
rect -3380 -14130 -3120 -14100
rect -3380 -14330 -3350 -14130
rect -3150 -14330 -3120 -14130
rect 11630 -14300 11660 -14100
rect 11860 -14300 11890 -14100
rect 11630 -14330 11890 -14300
rect -3380 -14360 -3120 -14330
rect 11630 -15130 11890 -15100
rect -3380 -15160 -3120 -15130
rect -3380 -15360 -3350 -15160
rect -3150 -15360 -3120 -15160
rect 11630 -15330 11660 -15130
rect 11860 -15330 11890 -15130
rect 11630 -15360 11890 -15330
rect -3380 -15390 -3120 -15360
rect 11630 -16160 11890 -16130
rect -3380 -16190 -3120 -16160
rect -3380 -16390 -3350 -16190
rect -3150 -16390 -3120 -16190
rect 11630 -16360 11660 -16160
rect 11860 -16360 11890 -16160
rect 11630 -16390 11890 -16360
rect -3380 -16420 -3120 -16390
rect 11630 -17190 11890 -17160
rect -3380 -17220 -3120 -17190
rect -3380 -17420 -3350 -17220
rect -3150 -17420 -3120 -17220
rect 11630 -17390 11660 -17190
rect 11860 -17390 11890 -17190
rect 11630 -17420 11890 -17390
rect -3380 -17450 -3120 -17420
rect 11630 -18220 11890 -18190
rect -3380 -18250 -3120 -18220
rect -3380 -18450 -3350 -18250
rect -3150 -18450 -3120 -18250
rect 11630 -18420 11660 -18220
rect 11860 -18420 11890 -18220
rect 11630 -18450 11890 -18420
rect -3380 -18480 -3120 -18450
rect 11630 -19250 11890 -19220
rect -3380 -19280 -3120 -19250
rect -3380 -19480 -3350 -19280
rect -3150 -19480 -3120 -19280
rect 11630 -19450 11660 -19250
rect 11860 -19450 11890 -19250
rect 11630 -19480 11890 -19450
rect -3380 -19510 -3120 -19480
rect -3380 -20430 -3120 -20400
rect -3380 -20630 -3350 -20430
rect -3150 -20630 -3120 -20430
rect -3380 -20660 -3120 -20630
rect -2480 -20430 -2220 -20400
rect -2480 -20630 -2450 -20430
rect -2250 -20630 -2220 -20430
rect -2480 -20660 -2220 -20630
rect -1450 -20430 -1190 -20400
rect -1450 -20630 -1420 -20430
rect -1220 -20630 -1190 -20430
rect -1450 -20660 -1190 -20630
rect -420 -20430 -160 -20400
rect -420 -20630 -390 -20430
rect -190 -20630 -160 -20430
rect -420 -20660 -160 -20630
rect 610 -20430 870 -20400
rect 610 -20630 640 -20430
rect 840 -20630 870 -20430
rect 610 -20660 870 -20630
rect 1640 -20430 1900 -20400
rect 1640 -20630 1670 -20430
rect 1870 -20630 1900 -20430
rect 1640 -20660 1900 -20630
rect 2670 -20430 2930 -20400
rect 2670 -20630 2700 -20430
rect 2900 -20630 2930 -20430
rect 2670 -20660 2930 -20630
rect 3700 -20430 3960 -20400
rect 3700 -20630 3730 -20430
rect 3930 -20630 3960 -20430
rect 3700 -20660 3960 -20630
rect 4730 -20430 4990 -20400
rect 4730 -20630 4760 -20430
rect 4960 -20630 4990 -20430
rect 4730 -20660 4990 -20630
rect 5760 -20430 6020 -20400
rect 5760 -20630 5790 -20430
rect 5990 -20630 6020 -20430
rect 5760 -20660 6020 -20630
rect 6790 -20430 7050 -20400
rect 6790 -20630 6820 -20430
rect 7020 -20630 7050 -20430
rect 6790 -20660 7050 -20630
rect 7820 -20430 8080 -20400
rect 7820 -20630 7850 -20430
rect 8050 -20630 8080 -20430
rect 7820 -20660 8080 -20630
rect 8850 -20430 9110 -20400
rect 8850 -20630 8880 -20430
rect 9080 -20630 9110 -20430
rect 8850 -20660 9110 -20630
rect 9880 -20430 10140 -20400
rect 9880 -20630 9910 -20430
rect 10110 -20630 10140 -20430
rect 9880 -20660 10140 -20630
rect 10910 -20430 11170 -20400
rect 10910 -20630 10940 -20430
rect 11140 -20630 11170 -20430
rect 10910 -20660 11170 -20630
rect 11630 -20430 11890 -20400
rect 11630 -20630 11660 -20430
rect 11860 -20630 11890 -20430
rect 11630 -20660 11890 -20630
<< psubdiffcont >>
rect -3350 330 -3150 530
rect -2450 330 -2250 530
rect -1420 330 -1220 530
rect -390 330 -190 530
rect 640 330 840 530
rect 1670 330 1870 530
rect 2700 330 2900 530
rect 3730 330 3930 530
rect 4760 330 4960 530
rect 5790 330 5990 530
rect 6820 330 7020 530
rect 7850 330 8050 530
rect 8880 330 9080 530
rect 9910 330 10110 530
rect 10940 330 11140 530
rect 11660 330 11860 530
rect -3350 -940 -3150 -740
rect 11660 -910 11860 -710
rect -3350 -1970 -3150 -1770
rect 11660 -1940 11860 -1740
rect -3350 -3000 -3150 -2800
rect -3350 -4030 -3150 -3830
rect -3350 -5060 -3150 -4860
rect 11660 -2970 11860 -2770
rect 11660 -4000 11860 -3800
rect 11660 -5030 11860 -4830
rect -3350 -6090 -3150 -5890
rect 11660 -6060 11860 -5860
rect -3350 -7120 -3150 -6920
rect 11660 -7090 11860 -6890
rect -3350 -8150 -3150 -7950
rect 11660 -8120 11860 -7920
rect -3350 -9180 -3150 -8980
rect 11660 -9150 11860 -8950
rect -3350 -10210 -3150 -10010
rect 11660 -10180 11860 -9980
rect -3350 -11240 -3150 -11040
rect 11660 -11210 11860 -11010
rect -3350 -12270 -3150 -12070
rect 11660 -12240 11860 -12040
rect -3350 -13300 -3150 -13100
rect 11660 -13270 11860 -13070
rect -3350 -14330 -3150 -14130
rect 11660 -14300 11860 -14100
rect -3350 -15360 -3150 -15160
rect 11660 -15330 11860 -15130
rect -3350 -16390 -3150 -16190
rect 11660 -16360 11860 -16160
rect -3350 -17420 -3150 -17220
rect 11660 -17390 11860 -17190
rect -3350 -18450 -3150 -18250
rect 11660 -18420 11860 -18220
rect -3350 -19480 -3150 -19280
rect 11660 -19450 11860 -19250
rect -3350 -20630 -3150 -20430
rect -2450 -20630 -2250 -20430
rect -1420 -20630 -1220 -20430
rect -390 -20630 -190 -20430
rect 640 -20630 840 -20430
rect 1670 -20630 1870 -20430
rect 2700 -20630 2900 -20430
rect 3730 -20630 3930 -20430
rect 4760 -20630 4960 -20430
rect 5790 -20630 5990 -20430
rect 6820 -20630 7020 -20430
rect 7850 -20630 8050 -20430
rect 8880 -20630 9080 -20430
rect 9910 -20630 10110 -20430
rect 10940 -20630 11140 -20430
rect 11660 -20630 11860 -20430
<< xpolycontact >>
rect 3976 -2998 4046 -2566
rect 3976 -5230 4046 -4798
rect 4294 -2998 4364 -2566
rect 4294 -5230 4364 -4798
<< xpolyres >>
rect 3976 -4798 4046 -2998
rect 4294 -4798 4364 -2998
<< locali >>
rect -3600 530 12130 780
rect -3600 330 -3350 530
rect -3150 330 -2450 530
rect -2250 330 -1420 530
rect -1220 330 -390 530
rect -190 330 640 530
rect 840 330 1670 530
rect 1870 330 2700 530
rect 2900 330 3730 530
rect 3930 330 4760 530
rect 4960 330 5790 530
rect 5990 330 6820 530
rect 7020 330 7850 530
rect 8050 330 8880 530
rect 9080 330 9910 530
rect 10110 330 10940 530
rect 11140 330 11660 530
rect 11860 330 12130 530
rect -3600 60 12130 330
rect -3600 -740 -2880 60
rect -3600 -940 -3350 -740
rect -3150 -940 -2880 -740
rect -3600 -1770 -2880 -940
rect -3600 -1970 -3350 -1770
rect -3150 -1970 -2880 -1770
rect -3600 -2800 -2880 -1970
rect 11410 -710 12130 60
rect 11410 -910 11660 -710
rect 11860 -910 12130 -710
rect 11410 -1740 12130 -910
rect 11410 -1940 11660 -1740
rect 11860 -1940 12130 -1740
rect 4100 -2180 4430 -2160
rect 4100 -2380 4210 -2180
rect 4410 -2380 4430 -2180
rect 4100 -2400 4430 -2380
rect -3600 -3000 -3350 -2800
rect -3150 -3000 -2880 -2800
rect 11410 -2770 12130 -1940
rect 11410 -2970 11660 -2770
rect 11860 -2970 12130 -2770
rect -3600 -3830 -2880 -3000
rect -3600 -4030 -3350 -3830
rect -3150 -4030 -2880 -3830
rect -3600 -4860 -2880 -4030
rect 11410 -3800 12130 -2970
rect 11410 -4000 11660 -3800
rect 11860 -4000 12130 -3800
rect -3600 -5060 -3350 -4860
rect -3150 -5060 -2880 -4860
rect -3600 -5890 -2880 -5060
rect 11410 -4830 12130 -4000
rect 11410 -5030 11660 -4830
rect 11860 -5030 12130 -4830
rect -3600 -6090 -3350 -5890
rect -3150 -6090 -2880 -5890
rect -3600 -6920 -2880 -6090
rect -3600 -7120 -3350 -6920
rect -3150 -7120 -2880 -6920
rect -3600 -7950 -2880 -7120
rect -3600 -8150 -3350 -7950
rect -3150 -8150 -2880 -7950
rect -3600 -8980 -2880 -8150
rect -3600 -9180 -3350 -8980
rect -3150 -9180 -2880 -8980
rect -3600 -10010 -2880 -9180
rect -3600 -10210 -3350 -10010
rect -3150 -10210 -2880 -10010
rect -3600 -11040 -2880 -10210
rect -3600 -11240 -3350 -11040
rect -3150 -11240 -2880 -11040
rect -3600 -12070 -2880 -11240
rect -3600 -12270 -3350 -12070
rect -3150 -12270 -2880 -12070
rect -3600 -13100 -2880 -12270
rect -3600 -13300 -3350 -13100
rect -3150 -13300 -2880 -13100
rect -3600 -14130 -2880 -13300
rect -3600 -14330 -3350 -14130
rect -3150 -14330 -2880 -14130
rect -3600 -15160 -2880 -14330
rect -3600 -15360 -3350 -15160
rect -3150 -15360 -2880 -15160
rect -3600 -16190 -2880 -15360
rect -3600 -16390 -3350 -16190
rect -3150 -16390 -2880 -16190
rect -3600 -17220 -2880 -16390
rect -3600 -17420 -3350 -17220
rect -3150 -17420 -2880 -17220
rect -3600 -18250 -2880 -17420
rect -3600 -18450 -3350 -18250
rect -3150 -18450 -2880 -18250
rect -3600 -19280 -2880 -18450
rect -3600 -19480 -3350 -19280
rect -3150 -19480 -2880 -19280
rect -3600 -20180 -2880 -19480
rect 11410 -5860 12130 -5030
rect 11410 -6060 11660 -5860
rect 11860 -6060 12130 -5860
rect 11410 -6890 12130 -6060
rect 11410 -7090 11660 -6890
rect 11860 -7090 12130 -6890
rect 11410 -7920 12130 -7090
rect 11410 -8120 11660 -7920
rect 11860 -8120 12130 -7920
rect 11410 -8950 12130 -8120
rect 11410 -9150 11660 -8950
rect 11860 -9150 12130 -8950
rect 11410 -9980 12130 -9150
rect 11410 -10180 11660 -9980
rect 11860 -10180 12130 -9980
rect 11410 -11010 12130 -10180
rect 11410 -11210 11660 -11010
rect 11860 -11210 12130 -11010
rect 11410 -12040 12130 -11210
rect 11410 -12240 11660 -12040
rect 11860 -12240 12130 -12040
rect 11410 -13070 12130 -12240
rect 11410 -13270 11660 -13070
rect 11860 -13270 12130 -13070
rect 11410 -14100 12130 -13270
rect 11410 -14300 11660 -14100
rect 11860 -14300 12130 -14100
rect 11410 -15130 12130 -14300
rect 11410 -15330 11660 -15130
rect 11860 -15330 12130 -15130
rect 11410 -16160 12130 -15330
rect 11410 -16360 11660 -16160
rect 11860 -16360 12130 -16160
rect 11410 -17190 12130 -16360
rect 11410 -17390 11660 -17190
rect 11860 -17390 12130 -17190
rect 11410 -18220 12130 -17390
rect 11410 -18420 11660 -18220
rect 11860 -18420 12130 -18220
rect 11410 -19250 12130 -18420
rect 11410 -19450 11660 -19250
rect 11860 -19450 12130 -19250
rect 11410 -20180 12130 -19450
rect -3600 -20430 12130 -20180
rect -3600 -20630 -3350 -20430
rect -3150 -20630 -2450 -20430
rect -2250 -20630 -1420 -20430
rect -1220 -20630 -390 -20430
rect -190 -20630 640 -20430
rect 840 -20630 1670 -20430
rect 1870 -20630 2700 -20430
rect 2900 -20630 3730 -20430
rect 3930 -20630 4760 -20430
rect 4960 -20630 5790 -20430
rect 5990 -20630 6820 -20430
rect 7020 -20630 7850 -20430
rect 8050 -20630 8880 -20430
rect 9080 -20630 9910 -20430
rect 10110 -20630 10940 -20430
rect 11140 -20630 11660 -20430
rect 11860 -20630 12130 -20430
rect -3600 -20900 12130 -20630
<< viali >>
rect 4210 -2380 4410 -2180
rect 3992 -2981 4030 -2584
rect 4310 -2981 4348 -2584
rect 3992 -5212 4030 -4815
rect 4310 -5212 4348 -4815
rect 4450 -5110 4610 -4950
rect 3730 -20630 3930 -20430
<< metal1 >>
rect 4180 -2180 4650 -2150
rect 4180 -2380 4210 -2180
rect 4410 -2380 4650 -2180
rect 4180 -2410 4650 -2380
rect 3986 -2580 4036 -2572
rect 4304 -2580 4354 -2572
rect 3986 -2584 4354 -2580
rect 3986 -2981 3992 -2584
rect 4030 -2981 4310 -2584
rect 4348 -2981 4354 -2584
rect 3986 -2990 4354 -2981
rect 3986 -2993 4036 -2990
rect 4304 -2993 4354 -2990
rect 3970 -4803 4000 -4800
rect 3970 -4810 4036 -4803
rect 3670 -4815 4036 -4810
rect 3670 -4950 3992 -4815
rect 3670 -5110 3710 -4950
rect 3870 -5110 3992 -4950
rect 3670 -5212 3992 -5110
rect 4030 -5212 4036 -4815
rect 3670 -5224 4036 -5212
rect 4304 -4810 4354 -4803
rect 4430 -4810 4650 -2410
rect 4304 -4815 4650 -4810
rect 4304 -5212 4310 -4815
rect 4348 -4950 4650 -4815
rect 4348 -5110 4450 -4950
rect 4610 -5110 4650 -4950
rect 4348 -5212 4650 -5110
rect 4304 -5224 4650 -5212
rect 3670 -5230 4000 -5224
rect 4340 -5230 4650 -5224
rect 3710 -20430 3950 -20410
rect 3710 -20630 3730 -20430
rect 3930 -20630 3950 -20430
rect 3710 -20650 3950 -20630
<< via1 >>
rect 3710 -5110 3870 -4950
rect 4450 -5110 4610 -4950
rect 3730 -20630 3930 -20430
<< metal2 >>
rect 3690 -4950 3890 -4930
rect 3690 -5110 3710 -4950
rect 3870 -5110 3890 -4950
rect 3690 -5130 3890 -5110
rect 4430 -4950 4630 -4930
rect 4430 -5110 4450 -4950
rect 4610 -5110 4630 -4950
rect 4430 -5130 4630 -5110
rect 3710 -20430 3950 -20410
rect 3710 -20630 3730 -20430
rect 3930 -20630 3950 -20430
rect 3710 -20650 3950 -20630
<< via2 >>
rect 3710 -5110 3870 -4950
rect 4450 -5110 4610 -4950
rect 3730 -20630 3930 -20430
<< metal3 >>
rect -2560 -6220 3600 -1030
rect 4610 -4930 10830 -970
rect 3690 -4950 3890 -4930
rect 3690 -5110 3710 -4950
rect 3870 -5110 3890 -4950
rect 3690 -5130 3890 -5110
rect 4430 -4950 10830 -4930
rect 4430 -5110 4450 -4950
rect 4610 -5110 10830 -4950
rect 4430 -5130 10830 -5110
rect 4610 -6220 10830 -5130
rect -2560 -7270 10830 -6220
rect -2560 -20010 10180 -7270
rect 140 -20020 920 -20010
rect 3710 -20410 3940 -20010
rect 3710 -20430 3950 -20410
rect 3710 -20630 3730 -20430
rect 3930 -20630 3950 -20430
rect 3710 -20650 3950 -20630
<< via3 >>
rect 3710 -5110 3870 -4950
rect 4450 -5110 4610 -4950
<< mimcap >>
rect -2460 -1170 3540 -1130
rect -2460 -7090 -2420 -1170
rect 3500 -7090 3540 -1170
rect -2460 -7130 3540 -7090
rect 4770 -1170 10770 -1130
rect 4770 -7090 4810 -1170
rect 10730 -7090 10770 -1170
rect 4770 -7130 10770 -7090
rect 4120 -7380 10120 -7340
rect -2460 -7560 3540 -7520
rect -2460 -13480 -2420 -7560
rect 3500 -13480 3540 -7560
rect 4120 -13300 4160 -7380
rect 10080 -13300 10120 -7380
rect 4120 -13340 10120 -13300
rect -2460 -13520 3540 -13480
rect 4120 -13770 10120 -13730
rect -2460 -13870 3540 -13830
rect -2460 -19790 -2420 -13870
rect 3500 -19790 3540 -13870
rect 4120 -19690 4160 -13770
rect 10080 -19690 10120 -13770
rect 4120 -19730 10120 -19690
rect -2460 -19830 3540 -19790
<< mimcapcontact >>
rect -2420 -7090 3500 -1170
rect 4810 -7090 10730 -1170
rect -2420 -13480 3500 -7560
rect 4160 -13300 10080 -7380
rect -2420 -19790 3500 -13870
rect 4160 -19690 10080 -13770
<< metal4 >>
rect -2421 -1170 140 -1169
rect 920 -1170 3501 -1169
rect -2421 -7090 -2420 -1170
rect 3500 -4810 3501 -1170
rect 4809 -1170 7370 -1169
rect 8150 -1170 10731 -1169
rect 4809 -4810 4810 -1170
rect 3500 -4930 3830 -4810
rect 4490 -4930 4810 -4810
rect 3500 -4950 3890 -4930
rect 3500 -5110 3710 -4950
rect 3870 -5110 3890 -4950
rect 3500 -5130 3890 -5110
rect 4430 -4950 4810 -4930
rect 4430 -5110 4450 -4950
rect 4610 -5110 4810 -4950
rect 4430 -5130 4810 -5110
rect 3500 -5230 3830 -5130
rect 4490 -5230 4810 -5130
rect 3500 -7090 3501 -5230
rect -2421 -7091 3501 -7090
rect 4809 -7090 4810 -5230
rect 10730 -7090 10731 -1170
rect 4809 -7091 7370 -7090
rect 8150 -7091 10731 -7090
rect 140 -7559 920 -7091
rect 4159 -7380 6720 -7379
rect 7500 -7380 10081 -7379
rect -2421 -7560 3501 -7559
rect -2421 -13480 -2420 -7560
rect 3500 -13480 3501 -7560
rect 4159 -13300 4160 -7380
rect 10080 -13300 10081 -7380
rect 4159 -13301 10081 -13300
rect -2421 -13481 3501 -13480
rect 140 -13869 920 -13481
rect 6720 -13769 7500 -13301
rect 4159 -13770 10081 -13769
rect -2421 -13870 3501 -13869
rect -2421 -19790 -2420 -13870
rect 3500 -16470 3501 -13870
rect 4159 -16470 4160 -13770
rect 3500 -17340 4160 -16470
rect 3500 -19790 3501 -17340
rect 4159 -19690 4160 -17340
rect 10080 -19690 10081 -13770
rect 4159 -19691 6720 -19690
rect 7510 -19691 10081 -19690
rect -2421 -19791 140 -19790
rect 920 -19791 3501 -19790
<< labels >>
rlabel locali 4310 -20570 4310 -20570 1 gnd
rlabel locali 4310 -20570 4310 -20570 1 gnd!
rlabel locali 4130 -2280 4130 -2280 1 v
<< end >>
