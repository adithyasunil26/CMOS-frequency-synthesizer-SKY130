magic
tech sky130A
magscale 1 2
timestamp 1640749174
<< locali >>
rect 2090 6970 2460 7390
use sky130_fd_pr__res_xhigh_po_0p35_6YXUWP  sky130_fd_pr__res_xhigh_po_0p35_6YXUWP_0
timestamp 1640749174
transform 1 0 2117 0 1 5962
box -37 -1432 37 1432
use sky130_fd_pr__res_xhigh_po_0p35_6YXUWP  sky130_fd_pr__res_xhigh_po_0p35_6YXUWP_1
timestamp 1640749174
transform 1 0 2437 0 1 5962
box -37 -1432 37 1432
use sky130_fd_pr__cap_mim_m3_1_C2TDQN  sky130_fd_pr__cap_mim_m3_1_C2TDQN_0
timestamp 1640749174
transform 1 0 2440 0 1 -153340
box -3150 -157500 3149 157500
<< end >>
