magic
tech sky130A
timestamp 1640863034
<< metal2 >>
rect 262 -400 318 240
rect 853 -400 909 240
rect 1444 -400 1500 240
rect 2035 -400 2091 240
rect 2626 -400 2682 240
rect 3217 -400 3273 240
rect 3808 -400 3864 240
rect 4399 -400 4455 240
rect 4990 -400 5046 240
rect 5581 -400 5637 240
rect 6172 -400 6228 240
rect 6763 -400 6819 240
rect 7354 -400 7410 240
rect 7945 -400 8001 240
rect 8536 -400 8592 240
rect 9127 -400 9183 240
rect 9718 -400 9774 240
rect 10309 -400 10365 240
rect 10900 -400 10956 240
rect 11491 -400 11547 240
rect 12082 -400 12138 240
rect 12673 -400 12729 240
rect 13264 -400 13320 240
rect 13855 -400 13911 240
rect 14446 -400 14502 240
rect 15037 -400 15093 240
rect 15628 -400 15684 240
rect 16219 -400 16275 240
rect 16810 -400 16866 240
rect 17401 -400 17457 240
rect 17992 -400 18048 240
rect 18583 -400 18639 240
rect 19174 -400 19230 240
rect 19765 -400 19821 240
rect 20356 -400 20412 240
rect 20947 -400 21003 240
rect 21538 -400 21594 240
rect 22129 -400 22185 240
rect 22720 -400 22776 240
rect 23311 -400 23367 240
rect 23902 -400 23958 240
rect 24493 -400 24549 240
rect 25084 -400 25140 240
rect 25675 -400 25731 240
rect 26266 -400 26322 240
rect 26857 -400 26913 240
rect 27448 -400 27504 240
rect 28039 -400 28095 240
rect 28630 -400 28686 240
rect 29221 -400 29277 240
rect 29812 -400 29868 240
rect 30403 -400 30459 240
rect 30994 -400 31050 240
rect 31585 -400 31641 240
rect 32176 -400 32232 240
rect 32767 -400 32823 240
rect 33358 -400 33414 240
rect 33949 -400 34005 240
rect 34540 -400 34596 240
rect 35131 -400 35187 240
rect 35722 -400 35778 240
rect 36313 -400 36369 240
rect 36904 -400 36960 240
rect 37495 -400 37551 240
rect 38086 -400 38142 240
rect 38677 -400 38733 240
rect 39268 -400 39324 240
rect 39859 -400 39915 240
rect 40450 -400 40506 240
rect 41041 -400 41097 240
rect 41632 -400 41688 240
rect 42223 -400 42279 240
rect 42814 -400 42870 240
rect 43405 -400 43461 240
rect 43996 -400 44052 240
rect 44587 -400 44643 240
rect 45178 -400 45234 240
rect 45769 -400 45825 240
rect 46360 -400 46416 240
rect 46951 -400 47007 240
rect 47542 -400 47598 240
rect 48133 -400 48189 240
rect 48724 -400 48780 240
rect 49315 -400 49371 240
rect 49906 -400 49962 240
rect 50497 -400 50553 240
rect 51088 -400 51144 240
rect 51679 -400 51735 240
rect 52270 -400 52326 240
rect 52861 -400 52917 240
rect 53452 -400 53508 240
rect 54043 -400 54099 240
rect 54634 -400 54690 240
rect 55225 -400 55281 240
rect 55816 -400 55872 240
rect 56407 -400 56463 240
rect 56998 -400 57054 240
rect 57589 -400 57645 240
rect 58180 -400 58236 240
rect 58771 -400 58827 240
rect 59362 -400 59418 240
rect 59953 -400 60009 240
rect 60544 -400 60600 240
rect 61135 -400 61191 240
rect 61726 -400 61782 240
rect 62317 -400 62373 240
rect 62908 -400 62964 240
rect 63499 -400 63555 240
rect 64090 -400 64146 240
rect 64681 -400 64737 240
rect 65272 -400 65328 240
rect 65863 -400 65919 240
rect 66454 -400 66510 240
rect 67045 -400 67101 240
rect 67636 -400 67692 240
rect 68227 -400 68283 240
rect 68818 -400 68874 240
rect 69409 -400 69465 240
rect 70000 -400 70056 240
rect 70591 -400 70647 240
rect 71182 -400 71238 240
rect 71773 -400 71829 240
rect 72364 -400 72420 240
rect 72955 -400 73011 240
rect 73546 -400 73602 240
rect 74137 -400 74193 240
rect 74728 -400 74784 240
rect 75319 -400 75375 240
rect 75910 -400 75966 240
rect 76501 -400 76557 240
rect 77092 -400 77148 240
rect 77683 -400 77739 240
rect 78274 -400 78330 240
rect 78865 -400 78921 240
rect 79456 -400 79512 240
rect 80047 -400 80103 240
rect 80638 -400 80694 240
rect 81229 -400 81285 240
rect 81820 -400 81876 240
rect 82411 -400 82467 240
rect 83002 -400 83058 240
rect 83593 -400 83649 240
rect 84184 -400 84240 240
rect 84775 -400 84831 240
rect 85366 -400 85422 240
rect 85957 -400 86013 240
rect 86548 -400 86604 240
rect 87139 -400 87195 240
rect 87730 -400 87786 240
rect 88321 -400 88377 240
rect 88912 -400 88968 240
rect 89503 -400 89559 240
rect 90094 -400 90150 240
rect 90685 -400 90741 240
rect 91276 -400 91332 240
rect 91867 -400 91923 240
rect 92458 -400 92514 240
rect 93049 -400 93105 240
rect 93640 -400 93696 240
rect 94231 -400 94287 240
rect 94822 -400 94878 240
rect 95413 -400 95469 240
rect 96004 -400 96060 240
rect 96595 -400 96651 240
rect 97186 -400 97242 240
rect 97777 -400 97833 240
rect 98368 -400 98424 240
rect 98959 -400 99015 240
rect 99550 -400 99606 240
rect 100141 -400 100197 240
rect 100732 -400 100788 240
rect 101323 -400 101379 240
rect 101914 -400 101970 240
rect 102505 -400 102561 240
rect 103096 -400 103152 240
rect 103687 -400 103743 240
rect 104278 -400 104334 240
rect 104869 -400 104925 240
rect 105460 -400 105516 240
rect 106051 -400 106107 240
rect 106642 -400 106698 240
rect 107233 -400 107289 240
rect 107824 -400 107880 240
rect 108415 -400 108471 240
rect 109006 -400 109062 240
rect 109597 -400 109653 240
rect 110188 -400 110244 240
rect 110779 -400 110835 240
rect 111370 -400 111426 240
rect 111961 -400 112017 240
rect 112552 -400 112608 240
rect 113143 -400 113199 240
rect 113734 -400 113790 240
rect 114325 -400 114381 240
rect 114916 -400 114972 240
rect 115507 -400 115563 240
rect 116098 -400 116154 240
rect 116689 -400 116745 240
rect 117280 -400 117336 240
rect 117871 -400 117927 240
rect 118462 -400 118518 240
rect 119053 -400 119109 240
rect 119644 -400 119700 240
rect 120235 -400 120291 240
rect 120826 -400 120882 240
rect 121417 -400 121473 240
rect 122008 -400 122064 240
rect 122599 -400 122655 240
rect 123190 -400 123246 240
rect 123781 -400 123837 240
rect 124372 -400 124428 240
rect 124963 -400 125019 240
rect 125554 -400 125610 240
rect 126145 -400 126201 240
rect 126736 -400 126792 240
rect 127327 -400 127383 240
rect 127918 -400 127974 240
rect 128509 -400 128565 240
rect 129100 -400 129156 240
rect 129691 -400 129747 240
rect 130282 -400 130338 240
rect 130873 -400 130929 240
rect 131464 -400 131520 240
rect 132055 -400 132111 240
rect 132646 -400 132702 240
rect 133237 -400 133293 240
rect 133828 -400 133884 240
rect 134419 -400 134475 240
rect 135010 -400 135066 240
rect 135601 -400 135657 240
rect 136192 -400 136248 240
rect 136783 -400 136839 240
rect 137374 -400 137430 240
rect 137965 -400 138021 240
rect 138556 -400 138612 240
rect 139147 -400 139203 240
rect 139738 -400 139794 240
rect 140329 -400 140385 240
rect 140920 -400 140976 240
rect 141511 -400 141567 240
rect 142102 -400 142158 240
rect 142693 -400 142749 240
rect 143284 -400 143340 240
rect 143875 -400 143931 240
rect 144466 -400 144522 240
rect 145057 -400 145113 240
rect 145648 -400 145704 240
rect 146239 -400 146295 240
rect 146830 -400 146886 240
rect 147421 -400 147477 240
rect 148012 -400 148068 240
rect 148603 -400 148659 240
rect 149194 -400 149250 240
rect 149785 -400 149841 240
rect 150376 -400 150432 240
rect 150967 -400 151023 240
rect 151558 -400 151614 240
rect 152149 -400 152205 240
rect 152740 -400 152796 240
rect 153331 -400 153387 240
rect 153922 -400 153978 240
rect 154513 -400 154569 240
rect 155104 -400 155160 240
rect 155695 -400 155751 240
rect 156286 -400 156342 240
rect 156877 -400 156933 240
rect 157468 -400 157524 240
rect 158059 -400 158115 240
rect 158650 -400 158706 240
rect 159241 -400 159297 240
rect 159832 -400 159888 240
rect 160423 -400 160479 240
rect 161014 -400 161070 240
rect 161605 -400 161661 240
rect 162196 -400 162252 240
rect 162787 -400 162843 240
rect 163378 -400 163434 240
rect 163969 -400 164025 240
rect 164560 -400 164616 240
rect 165151 -400 165207 240
rect 165742 -400 165798 240
rect 166333 -400 166389 240
rect 166924 -400 166980 240
rect 167515 -400 167571 240
rect 168106 -400 168162 240
rect 168697 -400 168753 240
rect 169288 -400 169344 240
rect 169879 -400 169935 240
rect 170470 -400 170526 240
rect 171061 -400 171117 240
rect 171652 -400 171708 240
rect 172243 -400 172299 240
rect 172834 -400 172890 240
rect 173425 -400 173481 240
rect 174016 -400 174072 240
rect 174607 -400 174663 240
rect 175198 -400 175254 240
rect 175789 -400 175845 240
rect 176380 -400 176436 240
rect 176971 -400 177027 240
rect 177562 -400 177618 240
rect 178153 -400 178209 240
rect 178744 -400 178800 240
rect 179335 -400 179391 240
rect 179926 -400 179982 240
rect 180517 -400 180573 240
rect 181108 -400 181164 240
rect 181699 -400 181755 240
rect 182290 -400 182346 240
rect 182881 -400 182937 240
rect 183472 -400 183528 240
rect 184063 -400 184119 240
rect 184654 -400 184710 240
rect 185245 -400 185301 240
rect 185836 -400 185892 240
rect 186427 -400 186483 240
rect 187018 -400 187074 240
rect 187609 -400 187665 240
rect 188200 -400 188256 240
rect 188791 -400 188847 240
rect 189382 -400 189438 240
rect 189973 -400 190029 240
rect 190564 -400 190620 240
rect 191155 -400 191211 240
rect 191746 -400 191802 240
rect 192337 -400 192393 240
rect 192928 -400 192984 240
rect 193519 -400 193575 240
rect 194110 -400 194166 240
rect 194701 -400 194757 240
rect 195292 -400 195348 240
rect 195883 -400 195939 240
rect 196474 -400 196530 240
rect 197065 -400 197121 240
rect 197656 -400 197712 240
rect 198247 -400 198303 240
rect 198838 -400 198894 240
rect 199429 -400 199485 240
rect 200020 -400 200076 240
rect 200611 -400 200667 240
rect 201202 -400 201258 240
rect 201793 -400 201849 240
rect 202384 -400 202440 240
rect 202975 -400 203031 240
rect 203566 -400 203622 240
rect 204157 -400 204213 240
rect 204748 -400 204804 240
rect 205339 -400 205395 240
rect 205930 -400 205986 240
rect 206521 -400 206577 240
rect 207112 -400 207168 240
rect 207703 -400 207759 240
rect 208294 -400 208350 240
rect 208885 -400 208941 240
rect 209476 -400 209532 240
rect 210067 -400 210123 240
rect 210658 -400 210714 240
rect 211249 -400 211305 240
rect 211840 -400 211896 240
rect 212431 -400 212487 240
rect 213022 -400 213078 240
rect 213613 -400 213669 240
rect 214204 -400 214260 240
rect 214795 -400 214851 240
rect 215386 -400 215442 240
rect 215977 -400 216033 240
rect 216568 -400 216624 240
rect 217159 -400 217215 240
rect 217750 -400 217806 240
rect 218341 -400 218397 240
rect 218932 -400 218988 240
rect 219523 -400 219579 240
rect 220114 -400 220170 240
rect 220705 -400 220761 240
rect 221296 -400 221352 240
rect 221887 -400 221943 240
rect 222478 -400 222534 240
rect 223069 -400 223125 240
rect 223660 -400 223716 240
rect 224251 -400 224307 240
rect 224842 -400 224898 240
rect 225433 -400 225489 240
rect 226024 -400 226080 240
rect 226615 -400 226671 240
rect 227206 -400 227262 240
rect 227797 -400 227853 240
rect 228388 -400 228444 240
rect 228979 -400 229035 240
rect 229570 -400 229626 240
rect 230161 -400 230217 240
rect 230752 -400 230808 240
rect 231343 -400 231399 240
rect 231934 -400 231990 240
rect 232525 -400 232581 240
rect 233116 -400 233172 240
rect 233707 -400 233763 240
rect 234298 -400 234354 240
rect 234889 -400 234945 240
rect 235480 -400 235536 240
rect 236071 -400 236127 240
rect 236662 -400 236718 240
rect 237253 -400 237309 240
rect 237844 -400 237900 240
rect 238435 -400 238491 240
rect 239026 -400 239082 240
rect 239617 -400 239673 240
rect 240208 -400 240264 240
rect 240799 -400 240855 240
rect 241390 -400 241446 240
rect 241981 -400 242037 240
rect 242572 -400 242628 240
rect 243163 -400 243219 240
rect 243754 -400 243810 240
rect 244345 -400 244401 240
rect 244936 -400 244992 240
rect 245527 -400 245583 240
rect 246118 -400 246174 240
rect 246709 -400 246765 240
rect 247300 -400 247356 240
rect 247891 -400 247947 240
rect 248482 -400 248538 240
rect 249073 -400 249129 240
rect 249664 -400 249720 240
rect 250255 -400 250311 240
rect 250846 -400 250902 240
rect 251437 -400 251493 240
rect 252028 -400 252084 240
rect 252619 -400 252675 240
rect 253210 -400 253266 240
rect 253801 -400 253857 240
rect 254392 -400 254448 240
rect 254983 -400 255039 240
rect 255574 -400 255630 240
rect 256165 -400 256221 240
rect 256756 -400 256812 240
rect 257347 -400 257403 240
rect 257938 -400 257994 240
rect 258529 -400 258585 240
rect 259120 -400 259176 240
rect 259711 -400 259767 240
rect 260302 -400 260358 240
rect 260893 -400 260949 240
rect 261484 -400 261540 240
rect 262075 -400 262131 240
rect 262666 -400 262722 240
rect 263257 -400 263313 240
rect 263848 -400 263904 240
rect 264439 -400 264495 240
rect 265030 -400 265086 240
rect 265621 -400 265677 240
rect 266212 -400 266268 240
rect 266803 -400 266859 240
rect 267394 -400 267450 240
rect 267985 -400 268041 240
rect 268576 -400 268632 240
rect 269167 -400 269223 240
rect 269758 -400 269814 240
rect 270349 -400 270405 240
rect 270940 -400 270996 240
rect 271531 -400 271587 240
rect 272122 -400 272178 240
rect 272713 -400 272769 240
rect 273304 -400 273360 240
rect 273895 -400 273951 240
rect 274486 -400 274542 240
rect 275077 -400 275133 240
rect 275668 -400 275724 240
rect 276259 -400 276315 240
rect 276850 -400 276906 240
rect 277441 -400 277497 240
rect 278032 -400 278088 240
rect 278623 -400 278679 240
rect 279214 -400 279270 240
rect 279805 -400 279861 240
rect 280396 -400 280452 240
rect 280987 -400 281043 240
rect 281578 -400 281634 240
rect 282169 -400 282225 240
rect 282760 -400 282816 240
rect 283351 -400 283407 240
rect 283942 -400 283998 240
rect 284533 -400 284589 240
rect 285124 -400 285180 240
rect 285715 -400 285771 240
rect 286306 -400 286362 240
rect 286897 -400 286953 240
rect 287488 -400 287544 240
rect 288079 -400 288135 240
rect 288670 -400 288726 240
rect 289261 -400 289317 240
rect 289852 -400 289908 240
rect 290443 -400 290499 240
rect 291034 -400 291090 240
rect 291625 -400 291681 240
<< metal3 >>
rect 8097 351150 10597 352400
rect 34097 351150 36597 352400
rect 60097 351150 62597 352400
rect 82797 351150 85297 352400
rect 85447 351150 86547 352400
rect 86697 351150 87797 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 111297 351150 112397 352400
rect 112547 351150 113647 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 162147 351150 163247 352400
rect 163397 351150 164497 352400
rect 164647 351150 167147 352400
rect 206697 351150 209197 352400
rect 232697 351150 235197 352400
rect 255297 351170 257697 352400
rect 260297 351170 262697 352400
rect 283297 351150 285797 352400
rect -400 340121 850 342621
rect 291150 338992 292400 341492
rect -400 321921 830 324321
rect 291170 319892 292400 322292
rect -400 316921 830 319321
rect 291170 314892 292400 317292
rect 291760 294736 292400 294792
rect 291760 294145 292400 294201
rect 291760 293554 292400 293610
rect 291760 292963 292400 293019
rect 291760 292372 292400 292428
rect 291760 291781 292400 291837
rect -400 279721 830 282121
rect -400 274721 830 277121
rect 291170 275281 292400 277681
rect 291170 270281 292400 272681
rect -400 255765 240 255821
rect -400 255174 240 255230
rect -400 254583 240 254639
rect -400 253992 240 254048
rect -400 253401 240 253457
rect -400 252810 240 252866
rect 291760 250025 292400 250081
rect 291760 249434 292400 249490
rect 291760 248843 292400 248899
rect 291760 248252 292400 248308
rect 291760 247661 292400 247717
rect 291760 247070 292400 247126
rect -400 234154 240 234210
rect -400 233563 240 233619
rect -400 232972 240 233028
rect -400 232381 240 232437
rect -400 231790 240 231846
rect -400 231199 240 231255
rect 291760 227814 292400 227870
rect 291760 227223 292400 227279
rect 291760 226632 292400 226688
rect 291760 226041 292400 226097
rect 291760 225450 292400 225506
rect 291760 224859 292400 224915
rect -400 212543 240 212599
rect -400 211952 240 212008
rect -400 211361 240 211417
rect -400 210770 240 210826
rect -400 210179 240 210235
rect -400 209588 240 209644
rect 291760 205603 292400 205659
rect 291760 205012 292400 205068
rect 291760 204421 292400 204477
rect 291760 203830 292400 203886
rect 291760 203239 292400 203295
rect 291760 202648 292400 202704
rect -400 190932 240 190988
rect -400 190341 240 190397
rect -400 189750 240 189806
rect -400 189159 240 189215
rect -400 188568 240 188624
rect -400 187977 240 188033
rect 291760 182392 292400 182448
rect 291760 181801 292400 181857
rect 291760 181210 292400 181266
rect 291760 180619 292400 180675
rect 291760 180028 292400 180084
rect 291760 179437 292400 179493
rect -400 169321 240 169377
rect -400 168730 240 168786
rect -400 168139 240 168195
rect -400 167548 240 167604
rect -400 166957 240 167013
rect -400 166366 240 166422
rect 291760 159781 292400 159837
rect 291760 159190 292400 159246
rect 291760 158599 292400 158655
rect 291760 158008 292400 158064
rect 291760 157417 292400 157473
rect 291760 156826 292400 156882
rect -400 147710 240 147766
rect -400 147119 240 147175
rect -400 146528 240 146584
rect -400 145937 240 145993
rect -400 145346 240 145402
rect -400 144755 240 144811
rect 291760 137570 292400 137626
rect 291760 136979 292400 137035
rect 291760 136388 292400 136444
rect 291760 135797 292400 135853
rect 291760 135206 292400 135262
rect 291760 134615 292400 134671
rect -400 126199 240 126255
rect -400 125608 240 125664
rect -400 125017 240 125073
rect -400 124426 240 124482
rect -400 123835 240 123891
rect -400 123244 240 123300
rect 291170 117615 292400 120015
rect 291170 112615 292400 115015
rect -400 107444 830 109844
rect -400 102444 830 104844
rect 291170 95715 292400 98115
rect 291170 90715 292400 93115
rect -400 86444 830 88844
rect -400 81444 830 83844
rect 291170 73415 292400 75815
rect 291170 68415 292400 70815
rect -400 62388 240 62444
rect -400 61797 240 61853
rect -400 61206 240 61262
rect -400 60615 240 60671
rect -400 60024 240 60080
rect -400 59433 240 59489
rect 291760 47559 292400 47615
rect 291760 46968 292400 47024
rect 291760 46377 292400 46433
rect 291760 45786 292400 45842
rect -400 40777 240 40833
rect -400 40186 240 40242
rect -400 39595 240 39651
rect -400 39004 240 39060
rect -400 38413 240 38469
rect -400 37822 240 37878
rect 291760 25230 292400 25286
rect 291760 24639 292400 24695
rect 291760 24048 292400 24104
rect 291760 23457 292400 23513
rect -400 19166 240 19222
rect -400 18575 240 18631
rect -400 17984 240 18040
rect -400 17393 240 17449
rect -400 16802 240 16858
rect -400 16211 240 16267
rect 291760 12001 292400 12057
rect 291760 11410 292400 11466
rect 291760 10819 292400 10875
rect 291760 10228 292400 10284
rect 291760 9637 292400 9693
rect 291760 9046 292400 9102
rect -400 8455 240 8511
rect 291760 8455 292400 8511
rect -400 7864 240 7920
rect 291760 7864 292400 7920
rect -400 7273 240 7329
rect 291760 7273 292400 7329
rect -400 6682 240 6738
rect 291760 6682 292400 6738
rect -400 6091 240 6147
rect 291760 6091 292400 6147
rect -400 5500 240 5556
rect 291760 5500 292400 5556
rect -400 4909 240 4965
rect 291760 4909 292400 4965
rect -400 4318 240 4374
rect 291760 4318 292400 4374
rect -400 3727 240 3783
rect 291760 3727 292400 3783
rect -400 3136 240 3192
rect 291760 3136 292400 3192
rect -400 2545 240 2601
rect 291760 2545 292400 2601
rect -400 1954 240 2010
rect 291760 1954 292400 2010
rect -400 1363 240 1419
rect 291760 1363 292400 1419
rect -400 772 240 828
rect 291760 772 292400 828
<< metal4 >>
rect 82797 351150 85297 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 164647 351150 167147 352400
<< metal5 >>
rect 82797 351150 85297 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 164647 351150 167147 352400
<< comment >>
rect -50 352000 292050 352050
rect -50 0 0 352000
rect 292000 0 292050 352000
rect -50 -50 292050 0
use pd  pd_0 ../avadhani
timestamp 1640777101
transform 1 0 46233 0 1 340608
box -115 -730 1470 690
use divider  divider_0 ../avadhani
timestamp 1640857911
transform 1 0 58605 0 1 340399
box -185 -70 4395 1990
use ro_complete  ro_complete_0
timestamp 1640809734
transform 1 0 7163 0 1 344610
box 362 -5330 4455 1180
use cp  cp_0
timestamp 1640602475
transform 1 0 33315 0 1 341930
box -245 -1715 4500 2030
<< labels >>
flabel metal3 s 291760 134615 292400 134671 0 FreeSans 560 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -400 190932 240 190988 0 FreeSans 560 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -400 169321 240 169377 0 FreeSans 560 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -400 147710 240 147766 0 FreeSans 560 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -400 126199 240 126255 0 FreeSans 560 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -400 62388 240 62444 0 FreeSans 560 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -400 40777 240 40833 0 FreeSans 560 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -400 19166 240 19222 0 FreeSans 560 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -400 8455 240 8511 0 FreeSans 560 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 291760 156826 292400 156882 0 FreeSans 560 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 291760 179437 292400 179493 0 FreeSans 560 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 291760 202648 292400 202704 0 FreeSans 560 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 291760 224859 292400 224915 0 FreeSans 560 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 291760 247070 292400 247126 0 FreeSans 560 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 291760 291781 292400 291837 0 FreeSans 560 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -400 255765 240 255821 0 FreeSans 560 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -400 234154 240 234210 0 FreeSans 560 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -400 212543 240 212599 0 FreeSans 560 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 291760 135206 292400 135262 0 FreeSans 560 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -400 190341 240 190397 0 FreeSans 560 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -400 168730 240 168786 0 FreeSans 560 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -400 147119 240 147175 0 FreeSans 560 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -400 125608 240 125664 0 FreeSans 560 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -400 61797 240 61853 0 FreeSans 560 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -400 40186 240 40242 0 FreeSans 560 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -400 18575 240 18631 0 FreeSans 560 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -400 7864 240 7920 0 FreeSans 560 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 291760 157417 292400 157473 0 FreeSans 560 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 291760 180028 292400 180084 0 FreeSans 560 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 291760 203239 292400 203295 0 FreeSans 560 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 291760 225450 292400 225506 0 FreeSans 560 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 291760 247661 292400 247717 0 FreeSans 560 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 291760 292372 292400 292428 0 FreeSans 560 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -400 255174 240 255230 0 FreeSans 560 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -400 233563 240 233619 0 FreeSans 560 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -400 211952 240 212008 0 FreeSans 560 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 291150 338992 292400 341492 0 FreeSans 560 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 340121 850 342621 0 FreeSans 560 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 283297 351150 285797 352400 0 FreeSans 960 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 232697 351150 235197 352400 0 FreeSans 960 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 206697 351150 209197 352400 0 FreeSans 960 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 60097 351150 62597 352400 0 FreeSans 960 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 34097 351150 36597 352400 0 FreeSans 960 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 8097 351150 10597 352400 0 FreeSans 960 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 163397 351150 164497 352400 0 FreeSans 960 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 112547 351150 113647 352400 0 FreeSans 960 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 86697 351150 87797 352400 0 FreeSans 960 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 162147 351150 163247 352400 0 FreeSans 960 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 111297 351150 112397 352400 0 FreeSans 960 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 85447 351150 86547 352400 0 FreeSans 960 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 291760 1363 292400 1419 0 FreeSans 560 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 291760 204421 292400 204477 0 FreeSans 560 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 291760 226632 292400 226688 0 FreeSans 560 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 291760 248843 292400 248899 0 FreeSans 560 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 291760 293554 292400 293610 0 FreeSans 560 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -400 253992 240 254048 0 FreeSans 560 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -400 232381 240 232437 0 FreeSans 560 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -400 210770 240 210826 0 FreeSans 560 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -400 189159 240 189215 0 FreeSans 560 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -400 167548 240 167604 0 FreeSans 560 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -400 145937 240 145993 0 FreeSans 560 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 291760 3727 292400 3783 0 FreeSans 560 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -400 124426 240 124482 0 FreeSans 560 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -400 60615 240 60671 0 FreeSans 560 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -400 39004 240 39060 0 FreeSans 560 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -400 17393 240 17449 0 FreeSans 560 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -400 6682 240 6738 0 FreeSans 560 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -400 4318 240 4374 0 FreeSans 560 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -400 1954 240 2010 0 FreeSans 560 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 291760 6091 292400 6147 0 FreeSans 560 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 291760 8455 292400 8511 0 FreeSans 560 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 291760 10819 292400 10875 0 FreeSans 560 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 291760 24048 292400 24104 0 FreeSans 560 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 291760 46377 292400 46433 0 FreeSans 560 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 291760 136388 292400 136444 0 FreeSans 560 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 291760 158599 292400 158655 0 FreeSans 560 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 291760 181210 292400 181266 0 FreeSans 560 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 291760 772 292400 828 0 FreeSans 560 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 291760 203830 292400 203886 0 FreeSans 560 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 291760 226041 292400 226097 0 FreeSans 560 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 291760 248252 292400 248308 0 FreeSans 560 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 291760 292963 292400 293019 0 FreeSans 560 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -400 254583 240 254639 0 FreeSans 560 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -400 232972 240 233028 0 FreeSans 560 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -400 211361 240 211417 0 FreeSans 560 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -400 189750 240 189806 0 FreeSans 560 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -400 168139 240 168195 0 FreeSans 560 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -400 146528 240 146584 0 FreeSans 560 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 291760 3136 292400 3192 0 FreeSans 560 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -400 125017 240 125073 0 FreeSans 560 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -400 61206 240 61262 0 FreeSans 560 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -400 39595 240 39651 0 FreeSans 560 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -400 17984 240 18040 0 FreeSans 560 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -400 7273 240 7329 0 FreeSans 560 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -400 4909 240 4965 0 FreeSans 560 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -400 2545 240 2601 0 FreeSans 560 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 291760 5500 292400 5556 0 FreeSans 560 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 291760 7864 292400 7920 0 FreeSans 560 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 291760 10228 292400 10284 0 FreeSans 560 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 291760 23457 292400 23513 0 FreeSans 560 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 291760 45786 292400 45842 0 FreeSans 560 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 291760 135797 292400 135853 0 FreeSans 560 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 291760 158008 292400 158064 0 FreeSans 560 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 291760 180619 292400 180675 0 FreeSans 560 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 291760 2545 292400 2601 0 FreeSans 560 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 291760 205603 292400 205659 0 FreeSans 560 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 291760 227814 292400 227870 0 FreeSans 560 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 291760 250025 292400 250081 0 FreeSans 560 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 291760 294736 292400 294792 0 FreeSans 560 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -400 252810 240 252866 0 FreeSans 560 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -400 231199 240 231255 0 FreeSans 560 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -400 209588 240 209644 0 FreeSans 560 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -400 187977 240 188033 0 FreeSans 560 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -400 166366 240 166422 0 FreeSans 560 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -400 144755 240 144811 0 FreeSans 560 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 291760 4909 292400 4965 0 FreeSans 560 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -400 123244 240 123300 0 FreeSans 560 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -400 59433 240 59489 0 FreeSans 560 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -400 37822 240 37878 0 FreeSans 560 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -400 16211 240 16267 0 FreeSans 560 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -400 5500 240 5556 0 FreeSans 560 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -400 3136 240 3192 0 FreeSans 560 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -400 772 240 828 0 FreeSans 560 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 291760 7273 292400 7329 0 FreeSans 560 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 291760 9637 292400 9693 0 FreeSans 560 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 291760 12001 292400 12057 0 FreeSans 560 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 291760 25230 292400 25286 0 FreeSans 560 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 291760 47559 292400 47615 0 FreeSans 560 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 291760 137570 292400 137626 0 FreeSans 560 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 291760 159781 292400 159837 0 FreeSans 560 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 291760 182392 292400 182448 0 FreeSans 560 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 291760 1954 292400 2010 0 FreeSans 560 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 291760 205012 292400 205068 0 FreeSans 560 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 291760 227223 292400 227279 0 FreeSans 560 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 291760 249434 292400 249490 0 FreeSans 560 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 291760 294145 292400 294201 0 FreeSans 560 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -400 253401 240 253457 0 FreeSans 560 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -400 231790 240 231846 0 FreeSans 560 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -400 210179 240 210235 0 FreeSans 560 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -400 188568 240 188624 0 FreeSans 560 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -400 166957 240 167013 0 FreeSans 560 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -400 145346 240 145402 0 FreeSans 560 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 291760 4318 292400 4374 0 FreeSans 560 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -400 123835 240 123891 0 FreeSans 560 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -400 60024 240 60080 0 FreeSans 560 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -400 38413 240 38469 0 FreeSans 560 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -400 16802 240 16858 0 FreeSans 560 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -400 6091 240 6147 0 FreeSans 560 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -400 3727 240 3783 0 FreeSans 560 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -400 1363 240 1419 0 FreeSans 560 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 291760 6682 292400 6738 0 FreeSans 560 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 291760 9046 292400 9102 0 FreeSans 560 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 291760 11410 292400 11466 0 FreeSans 560 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 291760 24639 292400 24695 0 FreeSans 560 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 291760 46968 292400 47024 0 FreeSans 560 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 291760 136979 292400 137035 0 FreeSans 560 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 291760 159190 292400 159246 0 FreeSans 560 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 291760 181801 292400 181857 0 FreeSans 560 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 62908 -400 62964 240 0 FreeSans 560 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 240208 -400 240264 240 0 FreeSans 560 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 241981 -400 242037 240 0 FreeSans 560 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 243754 -400 243810 240 0 FreeSans 560 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 245527 -400 245583 240 0 FreeSans 560 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 247300 -400 247356 240 0 FreeSans 560 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 249073 -400 249129 240 0 FreeSans 560 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 250846 -400 250902 240 0 FreeSans 560 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 252619 -400 252675 240 0 FreeSans 560 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 254392 -400 254448 240 0 FreeSans 560 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 256165 -400 256221 240 0 FreeSans 560 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 80638 -400 80694 240 0 FreeSans 560 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 257938 -400 257994 240 0 FreeSans 560 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 259711 -400 259767 240 0 FreeSans 560 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 261484 -400 261540 240 0 FreeSans 560 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 263257 -400 263313 240 0 FreeSans 560 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 265030 -400 265086 240 0 FreeSans 560 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 266803 -400 266859 240 0 FreeSans 560 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 268576 -400 268632 240 0 FreeSans 560 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 270349 -400 270405 240 0 FreeSans 560 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 272122 -400 272178 240 0 FreeSans 560 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 273895 -400 273951 240 0 FreeSans 560 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 82411 -400 82467 240 0 FreeSans 560 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 275668 -400 275724 240 0 FreeSans 560 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 277441 -400 277497 240 0 FreeSans 560 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 279214 -400 279270 240 0 FreeSans 560 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 280987 -400 281043 240 0 FreeSans 560 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 282760 -400 282816 240 0 FreeSans 560 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 284533 -400 284589 240 0 FreeSans 560 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 286306 -400 286362 240 0 FreeSans 560 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 288079 -400 288135 240 0 FreeSans 560 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 84184 -400 84240 240 0 FreeSans 560 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 85957 -400 86013 240 0 FreeSans 560 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 87730 -400 87786 240 0 FreeSans 560 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 89503 -400 89559 240 0 FreeSans 560 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 91276 -400 91332 240 0 FreeSans 560 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 93049 -400 93105 240 0 FreeSans 560 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 94822 -400 94878 240 0 FreeSans 560 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 96595 -400 96651 240 0 FreeSans 560 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 64681 -400 64737 240 0 FreeSans 560 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 98368 -400 98424 240 0 FreeSans 560 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 100141 -400 100197 240 0 FreeSans 560 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 101914 -400 101970 240 0 FreeSans 560 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 103687 -400 103743 240 0 FreeSans 560 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 105460 -400 105516 240 0 FreeSans 560 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 107233 -400 107289 240 0 FreeSans 560 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 109006 -400 109062 240 0 FreeSans 560 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 110779 -400 110835 240 0 FreeSans 560 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 112552 -400 112608 240 0 FreeSans 560 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 114325 -400 114381 240 0 FreeSans 560 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 66454 -400 66510 240 0 FreeSans 560 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 116098 -400 116154 240 0 FreeSans 560 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 117871 -400 117927 240 0 FreeSans 560 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 119644 -400 119700 240 0 FreeSans 560 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 121417 -400 121473 240 0 FreeSans 560 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 123190 -400 123246 240 0 FreeSans 560 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 124963 -400 125019 240 0 FreeSans 560 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 126736 -400 126792 240 0 FreeSans 560 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 128509 -400 128565 240 0 FreeSans 560 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 130282 -400 130338 240 0 FreeSans 560 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 132055 -400 132111 240 0 FreeSans 560 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 68227 -400 68283 240 0 FreeSans 560 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 133828 -400 133884 240 0 FreeSans 560 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 135601 -400 135657 240 0 FreeSans 560 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 137374 -400 137430 240 0 FreeSans 560 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 139147 -400 139203 240 0 FreeSans 560 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 140920 -400 140976 240 0 FreeSans 560 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 142693 -400 142749 240 0 FreeSans 560 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 144466 -400 144522 240 0 FreeSans 560 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 146239 -400 146295 240 0 FreeSans 560 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 148012 -400 148068 240 0 FreeSans 560 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 149785 -400 149841 240 0 FreeSans 560 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 70000 -400 70056 240 0 FreeSans 560 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 151558 -400 151614 240 0 FreeSans 560 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 153331 -400 153387 240 0 FreeSans 560 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 155104 -400 155160 240 0 FreeSans 560 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 156877 -400 156933 240 0 FreeSans 560 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 158650 -400 158706 240 0 FreeSans 560 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 160423 -400 160479 240 0 FreeSans 560 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 162196 -400 162252 240 0 FreeSans 560 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 163969 -400 164025 240 0 FreeSans 560 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 165742 -400 165798 240 0 FreeSans 560 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 167515 -400 167571 240 0 FreeSans 560 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 71773 -400 71829 240 0 FreeSans 560 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 169288 -400 169344 240 0 FreeSans 560 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 171061 -400 171117 240 0 FreeSans 560 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 172834 -400 172890 240 0 FreeSans 560 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 174607 -400 174663 240 0 FreeSans 560 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 176380 -400 176436 240 0 FreeSans 560 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 178153 -400 178209 240 0 FreeSans 560 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 179926 -400 179982 240 0 FreeSans 560 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 181699 -400 181755 240 0 FreeSans 560 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 183472 -400 183528 240 0 FreeSans 560 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 185245 -400 185301 240 0 FreeSans 560 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 73546 -400 73602 240 0 FreeSans 560 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 187018 -400 187074 240 0 FreeSans 560 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 188791 -400 188847 240 0 FreeSans 560 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 190564 -400 190620 240 0 FreeSans 560 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 192337 -400 192393 240 0 FreeSans 560 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 194110 -400 194166 240 0 FreeSans 560 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 195883 -400 195939 240 0 FreeSans 560 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 197656 -400 197712 240 0 FreeSans 560 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 199429 -400 199485 240 0 FreeSans 560 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 201202 -400 201258 240 0 FreeSans 560 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 202975 -400 203031 240 0 FreeSans 560 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 75319 -400 75375 240 0 FreeSans 560 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 204748 -400 204804 240 0 FreeSans 560 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 206521 -400 206577 240 0 FreeSans 560 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 208294 -400 208350 240 0 FreeSans 560 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 210067 -400 210123 240 0 FreeSans 560 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 211840 -400 211896 240 0 FreeSans 560 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 213613 -400 213669 240 0 FreeSans 560 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 215386 -400 215442 240 0 FreeSans 560 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 217159 -400 217215 240 0 FreeSans 560 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 218932 -400 218988 240 0 FreeSans 560 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 220705 -400 220761 240 0 FreeSans 560 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 77092 -400 77148 240 0 FreeSans 560 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 222478 -400 222534 240 0 FreeSans 560 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 224251 -400 224307 240 0 FreeSans 560 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 226024 -400 226080 240 0 FreeSans 560 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 227797 -400 227853 240 0 FreeSans 560 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 229570 -400 229626 240 0 FreeSans 560 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 231343 -400 231399 240 0 FreeSans 560 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 233116 -400 233172 240 0 FreeSans 560 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 234889 -400 234945 240 0 FreeSans 560 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 236662 -400 236718 240 0 FreeSans 560 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 238435 -400 238491 240 0 FreeSans 560 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 78865 -400 78921 240 0 FreeSans 560 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 63499 -400 63555 240 0 FreeSans 560 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 240799 -400 240855 240 0 FreeSans 560 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 242572 -400 242628 240 0 FreeSans 560 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 244345 -400 244401 240 0 FreeSans 560 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 246118 -400 246174 240 0 FreeSans 560 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 247891 -400 247947 240 0 FreeSans 560 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 249664 -400 249720 240 0 FreeSans 560 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 251437 -400 251493 240 0 FreeSans 560 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 253210 -400 253266 240 0 FreeSans 560 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 254983 -400 255039 240 0 FreeSans 560 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 256756 -400 256812 240 0 FreeSans 560 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 81229 -400 81285 240 0 FreeSans 560 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 258529 -400 258585 240 0 FreeSans 560 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 260302 -400 260358 240 0 FreeSans 560 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 262075 -400 262131 240 0 FreeSans 560 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 263848 -400 263904 240 0 FreeSans 560 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 265621 -400 265677 240 0 FreeSans 560 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 267394 -400 267450 240 0 FreeSans 560 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 269167 -400 269223 240 0 FreeSans 560 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 270940 -400 270996 240 0 FreeSans 560 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 272713 -400 272769 240 0 FreeSans 560 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 274486 -400 274542 240 0 FreeSans 560 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 83002 -400 83058 240 0 FreeSans 560 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 276259 -400 276315 240 0 FreeSans 560 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 278032 -400 278088 240 0 FreeSans 560 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 279805 -400 279861 240 0 FreeSans 560 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 281578 -400 281634 240 0 FreeSans 560 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 283351 -400 283407 240 0 FreeSans 560 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 285124 -400 285180 240 0 FreeSans 560 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 286897 -400 286953 240 0 FreeSans 560 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 288670 -400 288726 240 0 FreeSans 560 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 84775 -400 84831 240 0 FreeSans 560 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 86548 -400 86604 240 0 FreeSans 560 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 88321 -400 88377 240 0 FreeSans 560 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 90094 -400 90150 240 0 FreeSans 560 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 91867 -400 91923 240 0 FreeSans 560 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 93640 -400 93696 240 0 FreeSans 560 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 95413 -400 95469 240 0 FreeSans 560 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 97186 -400 97242 240 0 FreeSans 560 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 65272 -400 65328 240 0 FreeSans 560 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 98959 -400 99015 240 0 FreeSans 560 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 100732 -400 100788 240 0 FreeSans 560 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 102505 -400 102561 240 0 FreeSans 560 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 104278 -400 104334 240 0 FreeSans 560 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 106051 -400 106107 240 0 FreeSans 560 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 107824 -400 107880 240 0 FreeSans 560 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 109597 -400 109653 240 0 FreeSans 560 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 111370 -400 111426 240 0 FreeSans 560 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 113143 -400 113199 240 0 FreeSans 560 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 114916 -400 114972 240 0 FreeSans 560 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 67045 -400 67101 240 0 FreeSans 560 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 116689 -400 116745 240 0 FreeSans 560 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 118462 -400 118518 240 0 FreeSans 560 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 120235 -400 120291 240 0 FreeSans 560 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 122008 -400 122064 240 0 FreeSans 560 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 123781 -400 123837 240 0 FreeSans 560 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 125554 -400 125610 240 0 FreeSans 560 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 127327 -400 127383 240 0 FreeSans 560 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 129100 -400 129156 240 0 FreeSans 560 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 130873 -400 130929 240 0 FreeSans 560 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 132646 -400 132702 240 0 FreeSans 560 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 68818 -400 68874 240 0 FreeSans 560 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 134419 -400 134475 240 0 FreeSans 560 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 136192 -400 136248 240 0 FreeSans 560 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 137965 -400 138021 240 0 FreeSans 560 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 139738 -400 139794 240 0 FreeSans 560 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 141511 -400 141567 240 0 FreeSans 560 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 143284 -400 143340 240 0 FreeSans 560 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 145057 -400 145113 240 0 FreeSans 560 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 146830 -400 146886 240 0 FreeSans 560 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 148603 -400 148659 240 0 FreeSans 560 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 150376 -400 150432 240 0 FreeSans 560 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 70591 -400 70647 240 0 FreeSans 560 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 152149 -400 152205 240 0 FreeSans 560 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 153922 -400 153978 240 0 FreeSans 560 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 155695 -400 155751 240 0 FreeSans 560 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 157468 -400 157524 240 0 FreeSans 560 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 159241 -400 159297 240 0 FreeSans 560 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 161014 -400 161070 240 0 FreeSans 560 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 162787 -400 162843 240 0 FreeSans 560 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 164560 -400 164616 240 0 FreeSans 560 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 166333 -400 166389 240 0 FreeSans 560 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 168106 -400 168162 240 0 FreeSans 560 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 72364 -400 72420 240 0 FreeSans 560 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 169879 -400 169935 240 0 FreeSans 560 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 171652 -400 171708 240 0 FreeSans 560 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 173425 -400 173481 240 0 FreeSans 560 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 175198 -400 175254 240 0 FreeSans 560 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 176971 -400 177027 240 0 FreeSans 560 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 178744 -400 178800 240 0 FreeSans 560 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 180517 -400 180573 240 0 FreeSans 560 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 182290 -400 182346 240 0 FreeSans 560 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 184063 -400 184119 240 0 FreeSans 560 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 185836 -400 185892 240 0 FreeSans 560 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 74137 -400 74193 240 0 FreeSans 560 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 187609 -400 187665 240 0 FreeSans 560 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 189382 -400 189438 240 0 FreeSans 560 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 191155 -400 191211 240 0 FreeSans 560 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 192928 -400 192984 240 0 FreeSans 560 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 194701 -400 194757 240 0 FreeSans 560 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 196474 -400 196530 240 0 FreeSans 560 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 198247 -400 198303 240 0 FreeSans 560 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 200020 -400 200076 240 0 FreeSans 560 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 201793 -400 201849 240 0 FreeSans 560 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 203566 -400 203622 240 0 FreeSans 560 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 75910 -400 75966 240 0 FreeSans 560 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 205339 -400 205395 240 0 FreeSans 560 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 207112 -400 207168 240 0 FreeSans 560 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 208885 -400 208941 240 0 FreeSans 560 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 210658 -400 210714 240 0 FreeSans 560 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 212431 -400 212487 240 0 FreeSans 560 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 214204 -400 214260 240 0 FreeSans 560 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 215977 -400 216033 240 0 FreeSans 560 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 217750 -400 217806 240 0 FreeSans 560 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 219523 -400 219579 240 0 FreeSans 560 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 221296 -400 221352 240 0 FreeSans 560 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 77683 -400 77739 240 0 FreeSans 560 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 223069 -400 223125 240 0 FreeSans 560 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 224842 -400 224898 240 0 FreeSans 560 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 226615 -400 226671 240 0 FreeSans 560 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 228388 -400 228444 240 0 FreeSans 560 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 230161 -400 230217 240 0 FreeSans 560 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 231934 -400 231990 240 0 FreeSans 560 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 233707 -400 233763 240 0 FreeSans 560 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 235480 -400 235536 240 0 FreeSans 560 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 237253 -400 237309 240 0 FreeSans 560 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 239026 -400 239082 240 0 FreeSans 560 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 79456 -400 79512 240 0 FreeSans 560 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 64090 -400 64146 240 0 FreeSans 560 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 241390 -400 241446 240 0 FreeSans 560 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 243163 -400 243219 240 0 FreeSans 560 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 244936 -400 244992 240 0 FreeSans 560 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 246709 -400 246765 240 0 FreeSans 560 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 248482 -400 248538 240 0 FreeSans 560 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 250255 -400 250311 240 0 FreeSans 560 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 252028 -400 252084 240 0 FreeSans 560 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 253801 -400 253857 240 0 FreeSans 560 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 255574 -400 255630 240 0 FreeSans 560 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 257347 -400 257403 240 0 FreeSans 560 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 81820 -400 81876 240 0 FreeSans 560 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 259120 -400 259176 240 0 FreeSans 560 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 260893 -400 260949 240 0 FreeSans 560 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 262666 -400 262722 240 0 FreeSans 560 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 264439 -400 264495 240 0 FreeSans 560 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 266212 -400 266268 240 0 FreeSans 560 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 267985 -400 268041 240 0 FreeSans 560 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 269758 -400 269814 240 0 FreeSans 560 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 271531 -400 271587 240 0 FreeSans 560 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 273304 -400 273360 240 0 FreeSans 560 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 275077 -400 275133 240 0 FreeSans 560 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 83593 -400 83649 240 0 FreeSans 560 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 276850 -400 276906 240 0 FreeSans 560 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 278623 -400 278679 240 0 FreeSans 560 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 280396 -400 280452 240 0 FreeSans 560 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 282169 -400 282225 240 0 FreeSans 560 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 283942 -400 283998 240 0 FreeSans 560 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 285715 -400 285771 240 0 FreeSans 560 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 287488 -400 287544 240 0 FreeSans 560 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 289261 -400 289317 240 0 FreeSans 560 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 85366 -400 85422 240 0 FreeSans 560 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 87139 -400 87195 240 0 FreeSans 560 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 88912 -400 88968 240 0 FreeSans 560 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 90685 -400 90741 240 0 FreeSans 560 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 92458 -400 92514 240 0 FreeSans 560 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 94231 -400 94287 240 0 FreeSans 560 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 96004 -400 96060 240 0 FreeSans 560 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 97777 -400 97833 240 0 FreeSans 560 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 65863 -400 65919 240 0 FreeSans 560 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 99550 -400 99606 240 0 FreeSans 560 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 101323 -400 101379 240 0 FreeSans 560 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 103096 -400 103152 240 0 FreeSans 560 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 104869 -400 104925 240 0 FreeSans 560 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 106642 -400 106698 240 0 FreeSans 560 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 108415 -400 108471 240 0 FreeSans 560 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 110188 -400 110244 240 0 FreeSans 560 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 111961 -400 112017 240 0 FreeSans 560 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 113734 -400 113790 240 0 FreeSans 560 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 115507 -400 115563 240 0 FreeSans 560 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 67636 -400 67692 240 0 FreeSans 560 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 117280 -400 117336 240 0 FreeSans 560 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 119053 -400 119109 240 0 FreeSans 560 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 120826 -400 120882 240 0 FreeSans 560 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 122599 -400 122655 240 0 FreeSans 560 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 124372 -400 124428 240 0 FreeSans 560 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 126145 -400 126201 240 0 FreeSans 560 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 127918 -400 127974 240 0 FreeSans 560 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 129691 -400 129747 240 0 FreeSans 560 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 131464 -400 131520 240 0 FreeSans 560 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 133237 -400 133293 240 0 FreeSans 560 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 69409 -400 69465 240 0 FreeSans 560 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 135010 -400 135066 240 0 FreeSans 560 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 136783 -400 136839 240 0 FreeSans 560 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 138556 -400 138612 240 0 FreeSans 560 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 140329 -400 140385 240 0 FreeSans 560 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 142102 -400 142158 240 0 FreeSans 560 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 143875 -400 143931 240 0 FreeSans 560 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 145648 -400 145704 240 0 FreeSans 560 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 147421 -400 147477 240 0 FreeSans 560 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 149194 -400 149250 240 0 FreeSans 560 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 150967 -400 151023 240 0 FreeSans 560 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 71182 -400 71238 240 0 FreeSans 560 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 152740 -400 152796 240 0 FreeSans 560 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 154513 -400 154569 240 0 FreeSans 560 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 156286 -400 156342 240 0 FreeSans 560 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 158059 -400 158115 240 0 FreeSans 560 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 159832 -400 159888 240 0 FreeSans 560 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 161605 -400 161661 240 0 FreeSans 560 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 163378 -400 163434 240 0 FreeSans 560 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 165151 -400 165207 240 0 FreeSans 560 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 166924 -400 166980 240 0 FreeSans 560 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 168697 -400 168753 240 0 FreeSans 560 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 72955 -400 73011 240 0 FreeSans 560 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 170470 -400 170526 240 0 FreeSans 560 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 172243 -400 172299 240 0 FreeSans 560 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 174016 -400 174072 240 0 FreeSans 560 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 175789 -400 175845 240 0 FreeSans 560 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 177562 -400 177618 240 0 FreeSans 560 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 179335 -400 179391 240 0 FreeSans 560 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 181108 -400 181164 240 0 FreeSans 560 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 182881 -400 182937 240 0 FreeSans 560 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 184654 -400 184710 240 0 FreeSans 560 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 186427 -400 186483 240 0 FreeSans 560 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 74728 -400 74784 240 0 FreeSans 560 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 188200 -400 188256 240 0 FreeSans 560 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 189973 -400 190029 240 0 FreeSans 560 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 191746 -400 191802 240 0 FreeSans 560 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 193519 -400 193575 240 0 FreeSans 560 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 195292 -400 195348 240 0 FreeSans 560 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 197065 -400 197121 240 0 FreeSans 560 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 198838 -400 198894 240 0 FreeSans 560 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 200611 -400 200667 240 0 FreeSans 560 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 202384 -400 202440 240 0 FreeSans 560 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 204157 -400 204213 240 0 FreeSans 560 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 76501 -400 76557 240 0 FreeSans 560 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 205930 -400 205986 240 0 FreeSans 560 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 207703 -400 207759 240 0 FreeSans 560 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 209476 -400 209532 240 0 FreeSans 560 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 211249 -400 211305 240 0 FreeSans 560 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 213022 -400 213078 240 0 FreeSans 560 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 214795 -400 214851 240 0 FreeSans 560 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 216568 -400 216624 240 0 FreeSans 560 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 218341 -400 218397 240 0 FreeSans 560 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 220114 -400 220170 240 0 FreeSans 560 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 221887 -400 221943 240 0 FreeSans 560 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 78274 -400 78330 240 0 FreeSans 560 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 223660 -400 223716 240 0 FreeSans 560 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 225433 -400 225489 240 0 FreeSans 560 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 227206 -400 227262 240 0 FreeSans 560 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 228979 -400 229035 240 0 FreeSans 560 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 230752 -400 230808 240 0 FreeSans 560 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 232525 -400 232581 240 0 FreeSans 560 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 234298 -400 234354 240 0 FreeSans 560 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 236071 -400 236127 240 0 FreeSans 560 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 237844 -400 237900 240 0 FreeSans 560 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 239617 -400 239673 240 0 FreeSans 560 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 80047 -400 80103 240 0 FreeSans 560 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 289852 -400 289908 240 0 FreeSans 560 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 290443 -400 290499 240 0 FreeSans 560 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 291034 -400 291090 240 0 FreeSans 560 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 291625 -400 291681 240 0 FreeSans 560 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 291170 319892 292400 322292 0 FreeSans 560 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 291170 314892 292400 317292 0 FreeSans 560 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 321921 830 324321 0 FreeSans 560 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 316921 830 319321 0 FreeSans 560 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 291170 270281 292400 272681 0 FreeSans 560 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 291170 275281 292400 277681 0 FreeSans 560 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 291170 117615 292400 120015 0 FreeSans 560 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 291170 112615 292400 115015 0 FreeSans 560 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 102444 830 104844 0 FreeSans 560 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 107444 830 109844 0 FreeSans 560 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 260297 351170 262697 352400 0 FreeSans 960 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 255297 351170 257697 352400 0 FreeSans 960 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 291170 73415 292400 75815 0 FreeSans 560 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 291170 68415 292400 70815 0 FreeSans 560 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 279721 830 282121 0 FreeSans 560 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 274721 830 277121 0 FreeSans 560 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 291170 95715 292400 98115 0 FreeSans 560 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 291170 90715 292400 93115 0 FreeSans 560 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 86444 830 88844 0 FreeSans 560 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 81444 830 83844 0 FreeSans 560 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 262 -400 318 240 0 FreeSans 560 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 853 -400 909 240 0 FreeSans 560 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 1444 -400 1500 240 0 FreeSans 560 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 3808 -400 3864 240 0 FreeSans 560 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 23902 -400 23958 240 0 FreeSans 560 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 25675 -400 25731 240 0 FreeSans 560 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 27448 -400 27504 240 0 FreeSans 560 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 29221 -400 29277 240 0 FreeSans 560 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 30994 -400 31050 240 0 FreeSans 560 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 32767 -400 32823 240 0 FreeSans 560 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 34540 -400 34596 240 0 FreeSans 560 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 36313 -400 36369 240 0 FreeSans 560 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 38086 -400 38142 240 0 FreeSans 560 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 39859 -400 39915 240 0 FreeSans 560 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 6172 -400 6228 240 0 FreeSans 560 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 41632 -400 41688 240 0 FreeSans 560 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 43405 -400 43461 240 0 FreeSans 560 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 45178 -400 45234 240 0 FreeSans 560 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 46951 -400 47007 240 0 FreeSans 560 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 48724 -400 48780 240 0 FreeSans 560 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 50497 -400 50553 240 0 FreeSans 560 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 52270 -400 52326 240 0 FreeSans 560 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 54043 -400 54099 240 0 FreeSans 560 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 55816 -400 55872 240 0 FreeSans 560 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 57589 -400 57645 240 0 FreeSans 560 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 8536 -400 8592 240 0 FreeSans 560 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 59362 -400 59418 240 0 FreeSans 560 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 61135 -400 61191 240 0 FreeSans 560 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 10900 -400 10956 240 0 FreeSans 560 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 13264 -400 13320 240 0 FreeSans 560 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 15037 -400 15093 240 0 FreeSans 560 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 16810 -400 16866 240 0 FreeSans 560 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 18583 -400 18639 240 0 FreeSans 560 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 20356 -400 20412 240 0 FreeSans 560 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 22129 -400 22185 240 0 FreeSans 560 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 2035 -400 2091 240 0 FreeSans 560 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 4399 -400 4455 240 0 FreeSans 560 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 24493 -400 24549 240 0 FreeSans 560 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 26266 -400 26322 240 0 FreeSans 560 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 28039 -400 28095 240 0 FreeSans 560 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 29812 -400 29868 240 0 FreeSans 560 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 31585 -400 31641 240 0 FreeSans 560 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 33358 -400 33414 240 0 FreeSans 560 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 35131 -400 35187 240 0 FreeSans 560 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 36904 -400 36960 240 0 FreeSans 560 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 38677 -400 38733 240 0 FreeSans 560 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 40450 -400 40506 240 0 FreeSans 560 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 6763 -400 6819 240 0 FreeSans 560 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 42223 -400 42279 240 0 FreeSans 560 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 43996 -400 44052 240 0 FreeSans 560 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 45769 -400 45825 240 0 FreeSans 560 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 47542 -400 47598 240 0 FreeSans 560 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 49315 -400 49371 240 0 FreeSans 560 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 51088 -400 51144 240 0 FreeSans 560 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 52861 -400 52917 240 0 FreeSans 560 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 54634 -400 54690 240 0 FreeSans 560 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 56407 -400 56463 240 0 FreeSans 560 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 58180 -400 58236 240 0 FreeSans 560 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 9127 -400 9183 240 0 FreeSans 560 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 59953 -400 60009 240 0 FreeSans 560 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 61726 -400 61782 240 0 FreeSans 560 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 11491 -400 11547 240 0 FreeSans 560 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 13855 -400 13911 240 0 FreeSans 560 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 15628 -400 15684 240 0 FreeSans 560 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 17401 -400 17457 240 0 FreeSans 560 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 19174 -400 19230 240 0 FreeSans 560 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 20947 -400 21003 240 0 FreeSans 560 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 22720 -400 22776 240 0 FreeSans 560 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 4990 -400 5046 240 0 FreeSans 560 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 25084 -400 25140 240 0 FreeSans 560 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 26857 -400 26913 240 0 FreeSans 560 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 28630 -400 28686 240 0 FreeSans 560 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 30403 -400 30459 240 0 FreeSans 560 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 32176 -400 32232 240 0 FreeSans 560 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 33949 -400 34005 240 0 FreeSans 560 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 35722 -400 35778 240 0 FreeSans 560 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 37495 -400 37551 240 0 FreeSans 560 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 39268 -400 39324 240 0 FreeSans 560 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 41041 -400 41097 240 0 FreeSans 560 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 7354 -400 7410 240 0 FreeSans 560 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 42814 -400 42870 240 0 FreeSans 560 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 44587 -400 44643 240 0 FreeSans 560 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 46360 -400 46416 240 0 FreeSans 560 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 48133 -400 48189 240 0 FreeSans 560 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 49906 -400 49962 240 0 FreeSans 560 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 51679 -400 51735 240 0 FreeSans 560 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 53452 -400 53508 240 0 FreeSans 560 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 55225 -400 55281 240 0 FreeSans 560 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 56998 -400 57054 240 0 FreeSans 560 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 58771 -400 58827 240 0 FreeSans 560 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 9718 -400 9774 240 0 FreeSans 560 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 60544 -400 60600 240 0 FreeSans 560 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 62317 -400 62373 240 0 FreeSans 560 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 12082 -400 12138 240 0 FreeSans 560 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 14446 -400 14502 240 0 FreeSans 560 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 16219 -400 16275 240 0 FreeSans 560 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 17992 -400 18048 240 0 FreeSans 560 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 19765 -400 19821 240 0 FreeSans 560 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 21538 -400 21594 240 0 FreeSans 560 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 23311 -400 23367 240 0 FreeSans 560 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 5581 -400 5637 240 0 FreeSans 560 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 7945 -400 8001 240 0 FreeSans 560 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 10309 -400 10365 240 0 FreeSans 560 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 12673 -400 12729 240 0 FreeSans 560 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 2626 -400 2682 240 0 FreeSans 560 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 3217 -400 3273 240 0 FreeSans 560 90 0 0 wbs_we_i
port 677 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 292000 352000
<< end >>
