* SPICE3 file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
X0 pd_0/UP pd_0/tspc_r_0/Qbar1 GND gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X1 pd_0/tspc_r_0/Qbar pd_0/UP GND gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X2 pd_0/tspc_r_0/Z1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3 pd_0/UP pd_0/tspc_r_0/Qbar1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X4 pd_0/tspc_r_0/Qbar1 pd_0/REF pd_0/tspc_r_0/z5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X5 pd_0/tspc_r_0/z5 pd_0/tspc_r_0/Z3 GND gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X6 pd_0/tspc_r_0/Z3 pd_0/REF VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X7 pd_0/tspc_r_0/Z2 pd_0/REF pd_0/tspc_r_0/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X8 pd_0/tspc_r_0/Z3 pd_0/tspc_r_0/Z2 pd_0/tspc_r_0/Z4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X9 pd_0/tspc_r_0/Z4 pd_0/REF GND gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X10 pd_0/tspc_r_0/Z3 pd_0/R GND gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X11 pd_0/tspc_r_0/Qbar pd_0/UP VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X12 pd_0/tspc_r_0/Qbar1 pd_0/tspc_r_0/Z3 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X13 pd_0/tspc_r_0/Z2 VDD GND gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X14 pd_0/DOWN pd_0/tspc_r_1/Qbar1 GND gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X15 pd_0/tspc_r_1/Qbar pd_0/DOWN GND gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X16 pd_0/tspc_r_1/Z1 VDD VDD pd_0/tspc_r_1/w_n290_n40# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X17 pd_0/DOWN pd_0/tspc_r_1/Qbar1 VDD pd_0/tspc_r_1/w_n290_n40# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X18 pd_0/tspc_r_1/Qbar1 pd_0/DIV pd_0/tspc_r_1/z5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X19 pd_0/tspc_r_1/z5 pd_0/tspc_r_1/Z3 GND gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X20 pd_0/tspc_r_1/Z3 pd_0/DIV VDD pd_0/tspc_r_1/w_n290_n40# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X21 pd_0/tspc_r_1/Z2 pd_0/DIV pd_0/tspc_r_1/Z1 pd_0/tspc_r_1/w_n290_n40# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X22 pd_0/tspc_r_1/Z3 pd_0/tspc_r_1/Z2 pd_0/tspc_r_1/Z4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X23 pd_0/tspc_r_1/Z4 pd_0/DIV GND gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X24 pd_0/tspc_r_1/Z3 pd_0/R GND gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X25 pd_0/tspc_r_1/Qbar pd_0/DOWN VDD pd_0/tspc_r_1/w_n290_n40# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X26 pd_0/tspc_r_1/Qbar1 pd_0/tspc_r_1/Z3 VDD pd_0/tspc_r_1/w_n290_n40# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X27 pd_0/tspc_r_1/Z2 VDD GND gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X28 pd_0/R pd_0/and_pd_0/Out1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X29 pd_0/and_pd_0/Out1 pd_0/UP pd_0/and_pd_0/Z1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X30 pd_0/and_pd_0/Out1 pd_0/UP VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X31 pd_0/and_pd_0/Z1 pd_0/DOWN GND gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X32 pd_0/and_pd_0/Out1 pd_0/DOWN VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X33 pd_0/R pd_0/and_pd_0/Out1 GND gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X34 cp_0/a_7110_n2840# cp_0/down gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=1.8e+06u
X35 cp_0/a_7110_0# cp_0/upbar vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+07u l=1.8e+06u
X36 cp_0/a_10_n50# cp_0/vbias gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=1.8e+06u
X37 cp_0/a_10_n50# cp_0/a_10_n50# vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+07u l=1.8e+06u
X38 cp_0/a_3060_0# cp_0/a_1710_n2840# cp_0/a_1710_n2840# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+07u l=1.8e+06u
X39 vdd gnd cp_0/a_3060_0# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+07u l=1.8e+06u
X40 cp_0/a_3060_n2840# cp_0/a_1710_0# cp_0/a_1710_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=1.8e+06u
X41 cp_0/a_1710_n2840# cp_0/vbias gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=1.8e+06u
X42 gnd cp_0/out cp_0/a_3060_n2840# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=1.8e+06u
X43 cp_0/a_1710_0# cp_0/a_10_n50# vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+07u l=1.8e+06u
X44 cp_0/out cp_0/a_1710_n2840# cp_0/a_7110_0# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+07u l=1.8e+06u
X45 gnd vdd cp_0/a_3060_n2840# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=1.8e+06u
X46 cp_0/out cp_0/a_1710_0# cp_0/a_7110_n2840# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=9e+06u l=1.8e+06u
X47 vdd cp_0/out cp_0/a_3060_0# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+07u l=1.8e+06u
X48 ro_complete_0/cbank_0/v gnd gnd sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=1e+06u l=180000u
X49 ro_complete_0/cbank_2/v gnd gnd sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=1e+06u l=180000u
X50 ro_complete_0/cbank_1/v ro_complete_0/cbank_0/v ro_complete_0/ro_var_extend_0/vdd ro_complete_0/ro_var_extend_0/vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X51 ro_complete_0/cbank_2/v ro_complete_0/cbank_1/v ro_complete_0/ro_var_extend_0/vdd ro_complete_0/ro_var_extend_0/vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X52 ro_complete_0/cbank_0/v ro_complete_0/cbank_2/v ro_complete_0/ro_var_extend_0/vdd ro_complete_0/ro_var_extend_0/vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=300000u
X53 ro_complete_0/cbank_1/v gnd gnd sky130_fd_pr__cap_var_lvt pd=0u ps=0u ad=0p as=0p w=1e+06u l=180000u
X54 ro_complete_0/cbank_1/v ro_complete_0/cbank_0/v gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X55 ro_complete_0/cbank_0/v ro_complete_0/cbank_2/v gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X56 ro_complete_0/cbank_2/v ro_complete_0/cbank_1/v gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X57 gnd ro_complete_0/a0 ro_complete_0/cbank_0/switch_0/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X58 gnd ro_complete_0/a1 ro_complete_0/cbank_0/switch_1/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X59 gnd ro_complete_0/a3 ro_complete_0/cbank_0/switch_3/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X60 gnd ro_complete_0/a2 ro_complete_0/cbank_0/switch_2/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X61 gnd ro_complete_0/a4 ro_complete_0/cbank_0/switch_4/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X62 gnd ro_complete_0/a5 ro_complete_0/cbank_0/switch_5/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X63 ro_complete_0/cbank_0/v ro_complete_0/cbank_0/switch_3/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X64 ro_complete_0/cbank_0/v gnd sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5.2e+06u
X65 ro_complete_0/cbank_0/v ro_complete_0/cbank_0/switch_5/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X66 ro_complete_0/cbank_0/v ro_complete_0/cbank_0/switch_4/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X67 ro_complete_0/cbank_0/v ro_complete_0/cbank_0/switch_0/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X68 ro_complete_0/cbank_0/v ro_complete_0/cbank_0/switch_1/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X69 ro_complete_0/cbank_0/v ro_complete_0/cbank_0/switch_2/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X70 gnd ro_complete_0/a0 ro_complete_0/cbank_1/switch_0/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X71 gnd ro_complete_0/a1 ro_complete_0/cbank_1/switch_1/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X72 gnd ro_complete_0/a3 ro_complete_0/cbank_1/switch_3/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X73 gnd ro_complete_0/a2 ro_complete_0/cbank_1/switch_2/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X74 gnd ro_complete_0/a4 ro_complete_0/cbank_1/switch_4/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X75 gnd ro_complete_0/a5 ro_complete_0/cbank_1/switch_5/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X76 ro_complete_0/cbank_1/v ro_complete_0/cbank_1/switch_3/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X77 ro_complete_0/cbank_1/v gnd sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5.2e+06u
X78 ro_complete_0/cbank_1/v ro_complete_0/cbank_1/switch_5/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X79 ro_complete_0/cbank_1/v ro_complete_0/cbank_1/switch_4/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X80 ro_complete_0/cbank_1/v ro_complete_0/cbank_1/switch_0/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X81 ro_complete_0/cbank_1/v ro_complete_0/cbank_1/switch_1/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X82 ro_complete_0/cbank_1/v ro_complete_0/cbank_1/switch_2/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X83 gnd ro_complete_0/a0 ro_complete_0/cbank_2/switch_0/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X84 gnd ro_complete_0/a1 ro_complete_0/cbank_2/switch_1/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X85 gnd ro_complete_0/a3 ro_complete_0/cbank_2/switch_3/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X86 gnd ro_complete_0/a2 ro_complete_0/cbank_2/switch_2/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X87 gnd ro_complete_0/a4 ro_complete_0/cbank_2/switch_4/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X88 gnd ro_complete_0/a5 ro_complete_0/cbank_2/switch_5/vin gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=7.2e+06u l=350000u
X89 ro_complete_0/cbank_2/v ro_complete_0/cbank_2/switch_3/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X90 ro_complete_0/cbank_2/v gnd sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5.2e+06u
X91 ro_complete_0/cbank_2/v ro_complete_0/cbank_2/switch_5/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X92 ro_complete_0/cbank_2/v ro_complete_0/cbank_2/switch_4/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X93 ro_complete_0/cbank_2/v ro_complete_0/cbank_2/switch_0/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X94 ro_complete_0/cbank_2/v ro_complete_0/cbank_2/switch_1/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X95 ro_complete_0/cbank_2/v ro_complete_0/cbank_2/switch_2/vin sky130_fd_pr__cap_mim_m3_1 l=2.8e+06u w=2.8e+06u
X96 divider_0/and_0/A divider_0/nor_0/B divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X97 divider_0/and_0/A divider_0/nor_0/A divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X98 divider_0/nor_0/Z1 divider_0/nor_0/A divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=150000u
X99 divider_0/and_0/A divider_0/nor_0/B divider_0/nor_0/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=150000u
X100 divider_0/and_0/B divider_0/nor_1/B divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X101 divider_0/and_0/B divider_0/mc2 divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X102 divider_0/nor_1/Z1 divider_0/mc2 divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=150000u
X103 divider_0/and_0/B divider_0/nor_1/B divider_0/nor_1/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=150000u
X104 divider_0/prescaler_0/tspc_0/Z3 divider_0/prescaler_0/tspc_0/Z2 divider_0/prescaler_0/tspc_0/Z4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X105 divider_0/prescaler_0/tspc_0/Z4 divider_0/clk divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X106 divider_0/prescaler_0/tspc_0/Z1 divider_0/prescaler_0/tspc_0/D divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X107 divider_0/prescaler_0/tspc_0/Z2 divider_0/prescaler_0/tspc_0/D divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X108 divider_0/prescaler_0/Out divider_0/prescaler_0/tspc_0/a_740_n680# divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X109 divider_0/prescaler_0/tspc_0/a_740_n680# divider_0/prescaler_0/tspc_0/Z3 divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X110 divider_0/prescaler_0/tspc_0/Z2 divider_0/clk divider_0/prescaler_0/tspc_0/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X111 divider_0/prescaler_0/Out divider_0/prescaler_0/tspc_0/a_740_n680# divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X112 divider_0/prescaler_0/tspc_0/a_740_n680# divider_0/clk divider_0/prescaler_0/tspc_0/a_630_n680# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X113 divider_0/prescaler_0/tspc_0/a_630_n680# divider_0/prescaler_0/tspc_0/Z3 divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X114 divider_0/prescaler_0/tspc_0/Z3 divider_0/clk divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.9e+06u l=150000u
X115 divider_0/prescaler_0/tspc_1/Z3 divider_0/prescaler_0/tspc_1/Z2 divider_0/prescaler_0/tspc_1/Z4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X116 divider_0/prescaler_0/tspc_1/Z4 divider_0/clk divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X117 divider_0/prescaler_0/tspc_1/Z1 divider_0/prescaler_0/Out divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X118 divider_0/prescaler_0/tspc_1/Z2 divider_0/prescaler_0/Out divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X119 divider_0/prescaler_0/tspc_1/Q divider_0/prescaler_0/m1_2700_2190# divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X120 divider_0/prescaler_0/m1_2700_2190# divider_0/prescaler_0/tspc_1/Z3 divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X121 divider_0/prescaler_0/tspc_1/Z2 divider_0/clk divider_0/prescaler_0/tspc_1/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X122 divider_0/prescaler_0/tspc_1/Q divider_0/prescaler_0/m1_2700_2190# divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X123 divider_0/prescaler_0/m1_2700_2190# divider_0/clk divider_0/prescaler_0/tspc_1/a_630_n680# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X124 divider_0/prescaler_0/tspc_1/a_630_n680# divider_0/prescaler_0/tspc_1/Z3 divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X125 divider_0/prescaler_0/tspc_1/Z3 divider_0/clk divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.9e+06u l=150000u
X126 divider_0/prescaler_0/tspc_2/Z3 divider_0/prescaler_0/tspc_2/Z2 divider_0/prescaler_0/tspc_2/Z4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X127 divider_0/prescaler_0/tspc_2/Z4 divider_0/clk divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X128 divider_0/prescaler_0/tspc_2/Z1 divider_0/prescaler_0/tspc_2/D divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X129 divider_0/prescaler_0/tspc_2/Z2 divider_0/prescaler_0/tspc_2/D divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X130 divider_0/prescaler_0/tspc_2/Q divider_0/prescaler_0/tspc_2/a_740_n680# divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X131 divider_0/prescaler_0/tspc_2/a_740_n680# divider_0/prescaler_0/tspc_2/Z3 divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X132 divider_0/prescaler_0/tspc_2/Z2 divider_0/clk divider_0/prescaler_0/tspc_2/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X133 divider_0/prescaler_0/tspc_2/Q divider_0/prescaler_0/tspc_2/a_740_n680# divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X134 divider_0/prescaler_0/tspc_2/a_740_n680# divider_0/clk divider_0/prescaler_0/tspc_2/a_630_n680# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X135 divider_0/prescaler_0/tspc_2/a_630_n680# divider_0/prescaler_0/tspc_2/Z3 divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X136 divider_0/prescaler_0/tspc_2/Z3 divider_0/clk divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.9e+06u l=150000u
X137 divider_0/prescaler_0/tspc_0/D divider_0/prescaler_0/tspc_2/Q divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X138 divider_0/prescaler_0/tspc_0/D divider_0/prescaler_0/tspc_1/Q divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X139 divider_0/prescaler_0/nand_0/z1 divider_0/prescaler_0/tspc_2/Q divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X140 divider_0/prescaler_0/tspc_0/D divider_0/prescaler_0/tspc_1/Q divider_0/prescaler_0/nand_0/z1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X141 divider_0/prescaler_0/tspc_2/D divider_0/and_0/OUT divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X142 divider_0/prescaler_0/tspc_2/D divider_0/prescaler_0/m1_2700_2190# divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X143 divider_0/prescaler_0/nand_1/z1 divider_0/and_0/OUT divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X144 divider_0/prescaler_0/tspc_2/D divider_0/prescaler_0/m1_2700_2190# divider_0/prescaler_0/nand_1/z1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X145 divider_0/tspc_0/Z3 divider_0/tspc_0/Z2 divider_0/tspc_0/Z4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X146 divider_0/tspc_0/Z4 divider_0/prescaler_0/Out divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X147 divider_0/tspc_0/Z1 divider_0/nor_0/A divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X148 divider_0/tspc_0/Z2 divider_0/nor_0/A divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X149 divider_0/tspc_0/Q divider_0/nor_0/A divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X150 divider_0/nor_0/A divider_0/tspc_0/Z3 divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X151 divider_0/tspc_0/Z2 divider_0/prescaler_0/Out divider_0/tspc_0/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X152 divider_0/tspc_0/Q divider_0/nor_0/A divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X153 divider_0/nor_0/A divider_0/prescaler_0/Out divider_0/tspc_0/a_630_n680# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X154 divider_0/tspc_0/a_630_n680# divider_0/tspc_0/Z3 divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X155 divider_0/tspc_0/Z3 divider_0/prescaler_0/Out divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.9e+06u l=150000u
X156 divider_0/tspc_1/Z3 divider_0/tspc_1/Z2 divider_0/tspc_1/Z4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X157 divider_0/tspc_1/Z4 divider_0/tspc_0/Q divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X158 divider_0/tspc_1/Z1 divider_0/nor_0/B divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X159 divider_0/tspc_1/Z2 divider_0/nor_0/B divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X160 divider_0/tspc_1/Q divider_0/nor_0/B divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X161 divider_0/nor_0/B divider_0/tspc_1/Z3 divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X162 divider_0/tspc_1/Z2 divider_0/tspc_0/Q divider_0/tspc_1/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X163 divider_0/tspc_1/Q divider_0/nor_0/B divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X164 divider_0/nor_0/B divider_0/tspc_0/Q divider_0/tspc_1/a_630_n680# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X165 divider_0/tspc_1/a_630_n680# divider_0/tspc_1/Z3 divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X166 divider_0/tspc_1/Z3 divider_0/tspc_0/Q divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.9e+06u l=150000u
X167 divider_0/tspc_2/Z3 divider_0/tspc_2/Z2 divider_0/tspc_2/Z4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X168 divider_0/tspc_2/Z4 divider_0/tspc_1/Q divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X169 divider_0/tspc_2/Z1 divider_0/nor_1/B divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X170 divider_0/tspc_2/Z2 divider_0/nor_1/B divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X171 divider_0/Out divider_0/nor_1/B divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X172 divider_0/nor_1/B divider_0/tspc_2/Z3 divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X173 divider_0/tspc_2/Z2 divider_0/tspc_1/Q divider_0/tspc_2/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X174 divider_0/Out divider_0/nor_1/B divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X175 divider_0/nor_1/B divider_0/tspc_1/Q divider_0/tspc_2/a_630_n680# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X176 divider_0/tspc_2/a_630_n680# divider_0/tspc_2/Z3 divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X177 divider_0/tspc_2/Z3 divider_0/tspc_1/Q divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.9e+06u l=150000u
X178 divider_0/and_0/OUT divider_0/and_0/out1 divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.8e+06u l=150000u
X179 divider_0/and_0/Z1 divider_0/and_0/A divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X180 divider_0/and_0/out1 divider_0/and_0/A divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.6e+06u l=150000u
X181 divider_0/and_0/out1 divider_0/and_0/B divider_0/and_0/Z1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X182 divider_0/and_0/OUT divider_0/and_0/out1 divider_0/gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X183 divider_0/and_0/out1 divider_0/and_0/B divider_0/vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.6e+06u l=150000u
C0 divider_0/vdd divider_0/and_0/Z1 0.01fF
C1 divider_0/tspc_2/Z1 divider_0/tspc_2/Z2 1.07fF
C2 divider_0/tspc_1/Q divider_0/tspc_2/Z3 0.45fF
C3 divider_0/nor_1/B divider_0/Out 0.22fF
C4 pd_0/REF pd_0/tspc_r_0/Z1 0.17fF
C5 pd_0/tspc_r_0/Qbar1 pd_0/UP 0.11fF
C6 divider_0/nor_0/A divider_0/tspc_0/Z1 0.03fF
C7 divider_0/prescaler_0/tspc_0/a_740_n680# divider_0/prescaler_0/tspc_1/Z4 0.01fF
C8 divider_0/prescaler_0/Out divider_0/prescaler_0/tspc_1/Q 0.91fF
C9 divider_0/prescaler_0/tspc_0/Z3 divider_0/vdd 0.67fF
C10 divider_0/prescaler_0/tspc_0/Z2 divider_0/prescaler_0/tspc_0/a_630_n680# 0.01fF
C11 ro_complete_0/a4 ro_complete_0/cbank_2/switch_4/vin 0.09fF
C12 divider_0/tspc_1/Z1 divider_0/vdd 0.58fF
C13 pd_0/tspc_r_0/Z2 pd_0/R 0.21fF
C14 io_clamp_low[2] io_analog[6] 0.53fF
C15 divider_0/mc2 divider_0/nor_0/A 0.04fF
C16 divider_0/prescaler_0/tspc_0/Z3 divider_0/prescaler_0/tspc_0/Z1 0.06fF
C17 ro_complete_0/cbank_0/switch_3/vin ro_complete_0/cbank_0/switch_4/vin 0.20fF
C18 divider_0/nor_0/A divider_0/prescaler_0/tspc_1/Q 0.03fF
C19 divider_0/gnd divider_0/tspc_1/Q 0.33fF
C20 divider_0/prescaler_0/tspc_0/D divider_0/prescaler_0/tspc_2/Q 0.04fF
C21 divider_0/prescaler_0/tspc_0/a_740_n680# divider_0/vdd 0.52fF
C22 divider_0/nor_0/B divider_0/tspc_2/Z4 0.02fF
C23 pd_0/DOWN pd_0/and_pd_0/Z1 0.19fF
C24 ro_complete_0/a0 ro_complete_0/cbank_1/v 0.05fF
C25 divider_0/gnd divider_0/and_0/Z1 0.41fF
C26 divider_0/prescaler_0/tspc_1/Z3 divider_0/prescaler_0/tspc_1/a_630_n680# 0.05fF
C27 divider_0/prescaler_0/tspc_0/Z3 divider_0/gnd 0.27fF
C28 ro_complete_0/cbank_0/v ro_complete_0/cbank_1/v 0.04fF
C29 divider_0/tspc_0/Z1 divider_0/vdd 0.58fF
C30 divider_0/prescaler_0/tspc_1/Z4 divider_0/prescaler_0/tspc_1/Q 0.16fF
C31 divider_0/prescaler_0/tspc_2/Z1 divider_0/prescaler_0/tspc_2/Z2 1.07fF
C32 divider_0/tspc_2/Z3 divider_0/tspc_2/a_630_n680# 0.05fF
C33 cp_0/a_1710_0# cp_0/out 0.84fF
C34 divider_0/gnd divider_0/prescaler_0/tspc_0/a_740_n680# 0.22fF
C35 divider_0/mc2 divider_0/vdd 0.06fF
C36 divider_0/tspc_1/Z2 divider_0/tspc_1/a_630_n680# 0.01fF
C37 divider_0/prescaler_0/tspc_2/Z2 divider_0/prescaler_0/tspc_2/D 0.09fF
C38 divider_0/prescaler_0/tspc_1/Q divider_0/vdd 0.64fF
C39 cp_0/a_10_n50# cp_0/vbias 0.19fF
C40 pd_0/tspc_r_0/Qbar pd_0/and_pd_0/Z1 0.02fF
C41 pd_0/tspc_r_1/Z3 pd_0/tspc_r_1/z5 0.11fF
C42 ro_complete_0/cbank_0/switch_4/vin ro_complete_0/a3 0.13fF
C43 ro_complete_0/cbank_0/switch_3/vin ro_complete_0/cbank_0/v 1.30fF
C44 divider_0/gnd divider_0/tspc_2/a_630_n680# 0.61fF
C45 divider_0/vdd divider_0/tspc_2/Z2 0.36fF
C46 pd_0/and_pd_0/Out1 pd_0/and_pd_0/Z1 0.18fF
C47 ro_complete_0/cbank_0/switch_5/vin ro_complete_0/a4 0.12fF
C48 ro_complete_0/cbank_1/switch_4/vin ro_complete_0/cbank_1/switch_5/vin 0.19fF
C49 ro_complete_0/cbank_1/switch_2/vin ro_complete_0/a2 0.09fF
C50 divider_0/and_0/OUT divider_0/and_0/out1 0.31fF
C51 divider_0/tspc_1/Q divider_0/tspc_2/Z4 0.15fF
C52 divider_0/tspc_2/Z2 divider_0/tspc_2/Z3 0.16fF
C53 cp_0/a_1710_0# cp_0/a_10_n50# 0.04fF
C54 pd_0/tspc_r_0/Z3 pd_0/tspc_r_0/Z2 0.25fF
C55 divider_0/gnd divider_0/mc2 1.02fF
C56 divider_0/prescaler_0/Out divider_0/tspc_0/Z2 0.11fF
C57 divider_0/gnd divider_0/prescaler_0/tspc_1/Q 0.83fF
C58 divider_0/prescaler_0/tspc_0/Z4 divider_0/vdd 0.01fF
C59 divider_0/prescaler_0/tspc_2/Z2 divider_0/vdd 0.37fF
C60 GND pd_0/tspc_r_1/Qbar 0.14fF
C61 pd_0/DIV pd_0/tspc_r_1/Z3 0.65fF
C62 divider_0/prescaler_0/tspc_0/Z4 divider_0/prescaler_0/tspc_0/Z1 0.00fF
C63 ro_complete_0/cbank_1/switch_3/vin ro_complete_0/cbank_1/switch_2/vin 0.20fF
C64 divider_0/gnd divider_0/tspc_2/Z2 0.16fF
C65 divider_0/nor_0/A divider_0/tspc_0/Z2 0.23fF
C66 divider_0/prescaler_0/tspc_0/D divider_0/vdd 0.90fF
C67 divider_0/prescaler_0/Out divider_0/prescaler_0/m1_2700_2190# 0.11fF
C68 divider_0/prescaler_0/tspc_0/D divider_0/prescaler_0/tspc_0/Z1 0.03fF
C69 divider_0/tspc_1/Z2 divider_0/tspc_0/Q 0.14fF
C70 divider_0/tspc_1/Z3 divider_0/nor_0/B 0.38fF
C71 divider_0/and_0/OUT divider_0/clk 0.04fF
C72 divider_0/prescaler_0/tspc_0/Z4 divider_0/gnd 0.44fF
C73 divider_0/nor_0/A divider_0/prescaler_0/m1_2700_2190# 0.01fF
C74 divider_0/gnd divider_0/prescaler_0/tspc_2/Z2 0.16fF
C75 ro_complete_0/cbank_1/switch_5/vin ro_complete_0/a4 0.12fF
C76 divider_0/tspc_0/Z1 divider_0/tspc_0/Z3 0.06fF
C77 divider_0/prescaler_0/m1_2700_2190# divider_0/prescaler_0/tspc_2/D 0.16fF
C78 divider_0/prescaler_0/tspc_2/Z2 divider_0/prescaler_0/tspc_2/Z3 0.16fF
C79 divider_0/prescaler_0/tspc_1/a_630_n680# divider_0/prescaler_0/tspc_1/Q 0.04fF
C80 divider_0/tspc_2/Z4 divider_0/tspc_2/a_630_n680# 0.12fF
C81 divider_0/tspc_1/Z4 divider_0/tspc_1/a_630_n680# 0.12fF
C82 GND pd_0/tspc_r_0/z5 0.57fF
C83 divider_0/gnd divider_0/prescaler_0/tspc_0/D 0.05fF
C84 ro_complete_0/a4 ro_complete_0/cbank_2/v 0.05fF
C85 divider_0/vdd divider_0/tspc_0/Z2 0.37fF
C86 divider_0/prescaler_0/tspc_2/Q divider_0/prescaler_0/nand_0/z1 0.01fF
C87 divider_0/prescaler_0/tspc_1/Z3 divider_0/clk 0.45fF
C88 divider_0/and_0/out1 divider_0/and_0/Z1 0.36fF
C89 GND pd_0/and_pd_0/Z1 0.19fF
C90 pd_0/DOWN pd_0/tspc_r_1/z5 0.03fF
C91 pd_0/tspc_r_1/Z2 pd_0/R 0.21fF
C92 ro_complete_0/cbank_1/switch_3/vin ro_complete_0/a2 0.14fF
C93 divider_0/prescaler_0/m1_2700_2190# divider_0/prescaler_0/tspc_1/Z4 0.08fF
C94 divider_0/prescaler_0/tspc_0/Z2 divider_0/vdd 0.37fF
C95 divider_0/and_0/A divider_0/nor_0/B 0.26fF
C96 divider_0/vdd divider_0/Out 0.61fF
C97 divider_0/prescaler_0/tspc_0/Z1 divider_0/prescaler_0/tspc_0/Z2 1.07fF
C98 divider_0/tspc_0/a_630_n680# divider_0/nor_0/B 0.01fF
C99 divider_0/prescaler_0/m1_2700_2190# divider_0/vdd 0.59fF
C100 divider_0/tspc_2/Z2 divider_0/tspc_2/Z4 0.36fF
C101 divider_0/tspc_2/Z3 divider_0/Out 0.05fF
C102 pd_0/tspc_r_0/Qbar1 pd_0/tspc_r_0/Qbar 0.01fF
C103 pd_0/REF GND 0.04fF
C104 divider_0/gnd divider_0/tspc_0/Z2 0.16fF
C105 divider_0/tspc_1/Z3 divider_0/tspc_1/Q 0.05fF
C106 io_clamp_low[2] io_clamp_high[2] 0.53fF
C107 pd_0/tspc_r_1/Z3 pd_0/tspc_r_1/Qbar1 0.38fF
C108 io_clamp_high[1] io_analog[5] 0.53fF
C109 divider_0/gnd divider_0/prescaler_0/tspc_0/Z2 0.16fF
C110 divider_0/gnd divider_0/Out 0.29fF
C111 divider_0/prescaler_0/tspc_0/Z3 divider_0/clk 0.64fF
C112 divider_0/tspc_0/Q divider_0/tspc_1/Z4 0.15fF
C113 divider_0/gnd divider_0/prescaler_0/m1_2700_2190# 0.22fF
C114 ro_complete_0/cbank_1/switch_1/vin ro_complete_0/cbank_1/v 1.30fF
C115 divider_0/mc2 divider_0/and_0/out1 0.06fF
C116 divider_0/tspc_1/Z3 divider_0/tspc_1/Z1 0.06fF
C117 divider_0/prescaler_0/tspc_0/a_740_n680# divider_0/clk 0.14fF
C118 divider_0/nor_0/Z1 divider_0/vdd 0.75fF
C119 divider_0/nor_0/A divider_0/tspc_1/Z2 0.15fF
C120 ro_complete_0/cbank_1/switch_5/vin ro_complete_0/cbank_1/v 1.44fF
C121 divider_0/prescaler_0/m1_2700_2190# divider_0/prescaler_0/nand_1/z1 0.07fF
C122 divider_0/prescaler_0/tspc_2/Z2 divider_0/prescaler_0/tspc_2/Z4 0.36fF
C123 divider_0/nor_1/B divider_0/and_0/B 0.29fF
C124 ro_complete_0/cbank_1/v ro_complete_0/cbank_2/v 1.36fF
C125 divider_0/tspc_0/Z2 divider_0/tspc_0/Z3 0.16fF
C126 divider_0/vdd divider_0/prescaler_0/nand_0/z1 0.01fF
C127 pd_0/tspc_r_1/Z2 pd_0/tspc_r_1/Z4 0.14fF
C128 divider_0/gnd divider_0/nor_0/Z1 0.01fF
C129 ro_complete_0/cbank_0/switch_2/vin ro_complete_0/cbank_0/v 1.30fF
C130 ro_complete_0/a0 ro_complete_0/cbank_0/switch_0/vin 0.09fF
C131 divider_0/prescaler_0/tspc_1/Z1 divider_0/prescaler_0/tspc_1/Z3 0.06fF
C132 divider_0/prescaler_0/m1_2700_2190# divider_0/prescaler_0/tspc_1/a_630_n680# 0.19fF
C133 divider_0/prescaler_0/tspc_1/Q divider_0/clk 0.60fF
C134 ro_complete_0/cbank_0/v ro_complete_0/cbank_0/switch_0/vin 1.30fF
C135 divider_0/tspc_1/Z2 divider_0/vdd 0.36fF
C136 divider_0/nor_1/B divider_0/tspc_1/a_630_n680# 0.00fF
C137 pd_0/REF pd_0/tspc_r_0/z5 0.04fF
C138 pd_0/tspc_r_0/Z1 pd_0/tspc_r_0/Z2 0.71fF
C139 pd_0/tspc_r_0/Z3 pd_0/tspc_r_0/Z4 0.20fF
C140 pd_0/tspc_r_0/Qbar1 GND 0.16fF
C141 divider_0/mc2 divider_0/prescaler_0/tspc_2/a_630_n680# 0.19fF
C142 divider_0/gnd divider_0/prescaler_0/nand_0/z1 0.16fF
C143 ro_complete_0/cbank_1/v ro_complete_0/a5 0.08fF
C144 ro_complete_0/cbank_2/switch_4/vin ro_complete_0/cbank_2/switch_5/vin 0.19fF
C145 divider_0/nor_1/Z1 divider_0/and_0/B 0.78fF
C146 pd_0/tspc_r_0/Z4 pd_0/tspc_r_1/Z4 0.02fF
C147 GND pd_0/tspc_r_1/z5 0.57fF
C148 pd_0/DIV pd_0/tspc_r_1/Z1 0.17fF
C149 pd_0/tspc_r_1/Qbar1 pd_0/DOWN 0.11fF
C150 io_clamp_low[0] io_analog[4] 0.53fF
C151 ro_complete_0/cbank_1/switch_3/vin ro_complete_0/cbank_1/switch_4/vin 0.20fF
C152 divider_0/prescaler_0/tspc_0/Z4 divider_0/clk 0.12fF
C153 divider_0/tspc_0/Q divider_0/tspc_1/a_630_n680# 0.01fF
C154 divider_0/prescaler_0/tspc_2/Z2 divider_0/clk 0.11fF
C155 divider_0/mc2 divider_0/and_0/A 0.16fF
C156 divider_0/gnd divider_0/tspc_1/Z2 0.16fF
C157 divider_0/nor_0/A divider_0/tspc_1/Z4 0.02fF
C158 divider_0/prescaler_0/tspc_0/D divider_0/clk 0.29fF
C159 ro_complete_0/a3 ro_complete_0/cbank_2/v 0.05fF
C160 divider_0/prescaler_0/tspc_2/a_740_n680# divider_0/prescaler_0/tspc_2/Q 0.20fF
C161 divider_0/prescaler_0/tspc_2/Z2 divider_0/prescaler_0/tspc_2/a_630_n680# 0.01fF
C162 GND pd_0/DIV 0.04fF
C163 pd_0/tspc_r_0/Z3 pd_0/R 0.35fF
C164 divider_0/nor_0/B divider_0/tspc_1/Q 0.51fF
C165 ro_complete_0/a3 ro_complete_0/cbank_2/switch_3/vin 0.09fF
C166 divider_0/vdd divider_0/tspc_1/Z4 0.01fF
C167 ro_complete_0/cbank_1/switch_2/vin ro_complete_0/cbank_1/v 1.30fF
C168 divider_0/nor_0/A divider_0/and_0/B 0.08fF
C169 divider_0/nor_0/B divider_0/tspc_1/Z1 0.03fF
C170 divider_0/prescaler_0/tspc_0/Z2 divider_0/clk 0.11fF
C171 divider_0/nor_1/Z1 divider_0/nor_1/B 0.06fF
C172 divider_0/and_0/OUT divider_0/and_0/Z1 0.04fF
C173 pd_0/tspc_r_0/Qbar1 pd_0/tspc_r_0/z5 0.20fF
C174 divider_0/prescaler_0/Out divider_0/tspc_0/Z4 0.12fF
C175 ro_complete_0/a1 ro_complete_0/cbank_2/v 0.05fF
C176 divider_0/prescaler_0/m1_2700_2190# divider_0/clk 0.01fF
C177 io_clamp_low[1] io_clamp_high[1] 0.53fF
C178 pd_0/tspc_r_0/z5 pd_0/tspc_r_1/z5 0.02fF
C179 pd_0/tspc_r_1/Z3 pd_0/tspc_r_1/Z2 0.25fF
C180 divider_0/gnd divider_0/tspc_1/Z4 0.44fF
C181 divider_0/nor_0/A divider_0/tspc_0/Z4 0.21fF
C182 divider_0/prescaler_0/Out divider_0/prescaler_0/tspc_1/Z2 0.19fF
C183 divider_0/nor_1/B divider_0/tspc_2/Z1 0.03fF
C184 divider_0/vdd divider_0/and_0/B 0.20fF
C185 cp_0/upbar cp_0/a_1710_n2840# 0.29fF
C186 pd_0/REF pd_0/tspc_r_0/Qbar1 0.12fF
C187 divider_0/mc2 divider_0/nor_0/B 0.07fF
C188 ro_complete_0/a2 ro_complete_0/cbank_1/v 0.05fF
C189 divider_0/tspc_0/a_630_n680# divider_0/tspc_0/Z2 0.01fF
C190 divider_0/prescaler_0/tspc_2/a_740_n680# divider_0/vdd 0.52fF
C191 cp_0/a_1710_0# cp_0/down 0.32fF
C192 pd_0/UP pd_0/R 0.45fF
C193 GND pd_0/tspc_r_1/Qbar1 0.16fF
C194 divider_0/mc2 divider_0/and_0/OUT 0.05fF
C195 ro_complete_0/cbank_2/switch_5/vin ro_complete_0/cbank_2/v 1.45fF
C196 divider_0/nor_0/B divider_0/tspc_2/Z2 0.20fF
C197 divider_0/vdd divider_0/tspc_0/Z4 0.01fF
C198 divider_0/prescaler_0/Out divider_0/prescaler_0/tspc_0/a_630_n680# 0.04fF
C199 ro_complete_0/cbank_0/switch_3/vin ro_complete_0/a2 0.14fF
C200 ro_complete_0/cbank_1/switch_3/vin ro_complete_0/cbank_1/v 1.30fF
C201 ro_complete_0/cbank_0/switch_4/vin ro_complete_0/cbank_0/v 1.30fF
C202 divider_0/prescaler_0/tspc_1/Z2 divider_0/prescaler_0/tspc_1/Z4 0.36fF
C203 divider_0/gnd divider_0/and_0/B 0.45fF
C204 divider_0/gnd divider_0/prescaler_0/tspc_2/a_740_n680# 0.22fF
C205 ro_complete_0/a0 ro_complete_0/cbank_2/switch_0/vin 0.09fF
C206 ro_complete_0/cbank_1/switch_4/vin ro_complete_0/a4 0.09fF
C207 divider_0/prescaler_0/tspc_2/a_740_n680# divider_0/prescaler_0/tspc_2/Z3 0.33fF
C208 divider_0/prescaler_0/tspc_1/Z2 divider_0/vdd 0.38fF
C209 divider_0/prescaler_0/tspc_1/Z3 divider_0/prescaler_0/tspc_1/Q 0.21fF
C210 divider_0/tspc_1/Q divider_0/tspc_2/a_630_n680# 0.01fF
C211 pd_0/tspc_r_0/Z2 GND 0.14fF
C212 divider_0/prescaler_0/tspc_0/Z3 divider_0/prescaler_0/tspc_0/a_740_n680# 0.33fF
C213 divider_0/nor_0/A divider_0/tspc_0/Q 0.55fF
C214 divider_0/gnd divider_0/tspc_0/Z4 0.44fF
C215 divider_0/nor_0/Z1 divider_0/and_0/A 0.80fF
C216 ro_complete_0/a5 ro_complete_0/cbank_2/switch_5/vin 0.09fF
C217 ro_complete_0/cbank_1/v ro_complete_0/cbank_1/switch_0/vin 1.30fF
C218 divider_0/prescaler_0/tspc_2/Z2 divider_0/and_0/OUT 0.05fF
C219 pd_0/tspc_r_1/Qbar1 pd_0/tspc_r_1/Qbar 0.01fF
C220 pd_0/tspc_r_1/Z3 pd_0/R 0.29fF
C221 divider_0/tspc_1/Z2 divider_0/tspc_1/Z3 0.16fF
C222 divider_0/gnd divider_0/tspc_1/a_630_n680# 0.62fF
C223 divider_0/vdd divider_0/nor_1/B 0.55fF
C224 divider_0/gnd divider_0/prescaler_0/tspc_1/Z2 0.17fF
C225 ro_complete_0/cbank_1/switch_2/vin ro_complete_0/a1 0.14fF
C226 divider_0/mc2 divider_0/and_0/Z1 0.09fF
C227 divider_0/tspc_1/Q divider_0/tspc_2/Z2 0.14fF
C228 divider_0/nor_1/B divider_0/tspc_2/Z3 0.38fF
C229 pd_0/tspc_r_0/Z3 pd_0/UP 0.03fF
C230 divider_0/prescaler_0/tspc_0/Z3 divider_0/prescaler_0/tspc_1/Q 0.13fF
C231 divider_0/tspc_0/Q divider_0/vdd 0.72fF
C232 ro_complete_0/cbank_1/switch_3/vin ro_complete_0/a3 0.09fF
C233 divider_0/prescaler_0/tspc_0/a_740_n680# divider_0/prescaler_0/tspc_1/Q 0.15fF
C234 divider_0/gnd divider_0/nor_1/B 0.96fF
C235 divider_0/tspc_0/Z3 divider_0/tspc_0/Z4 0.65fF
C236 divider_0/gnd divider_0/prescaler_0/tspc_0/a_630_n680# 0.63fF
C237 divider_0/prescaler_0/tspc_0/Z2 divider_0/and_0/OUT 0.06fF
C238 divider_0/prescaler_0/tspc_1/Z2 divider_0/prescaler_0/tspc_1/a_630_n680# 0.01fF
C239 divider_0/nor_1/Z1 divider_0/vdd 0.75fF
C240 divider_0/prescaler_0/tspc_0/Z3 divider_0/prescaler_0/tspc_0/Z4 0.65fF
C241 divider_0/gnd divider_0/tspc_0/Q 0.33fF
C242 ro_complete_0/cbank_1/switch_4/vin ro_complete_0/cbank_1/v 1.30fF
C243 divider_0/prescaler_0/m1_2700_2190# divider_0/and_0/OUT 0.14fF
C244 divider_0/prescaler_0/tspc_2/a_740_n680# divider_0/prescaler_0/tspc_2/Z4 0.08fF
C245 divider_0/tspc_2/Z2 divider_0/tspc_2/a_630_n680# 0.01fF
C246 divider_0/prescaler_0/Out divider_0/nor_0/A 0.15fF
C247 divider_0/prescaler_0/tspc_0/Z3 divider_0/prescaler_0/tspc_0/D 0.05fF
C248 divider_0/prescaler_0/tspc_0/Z4 divider_0/prescaler_0/tspc_0/a_740_n680# 0.08fF
C249 ro_complete_0/cbank_2/switch_2/vin ro_complete_0/cbank_2/v 1.30fF
C250 divider_0/tspc_1/Z3 divider_0/tspc_1/Z4 0.65fF
C251 divider_0/prescaler_0/tspc_2/Q divider_0/vdd 0.70fF
C252 divider_0/prescaler_0/tspc_2/Z1 divider_0/prescaler_0/tspc_2/D 0.15fF
C253 divider_0/and_0/out1 divider_0/and_0/B 0.18fF
C254 io_clamp_low[0] io_clamp_high[0] 0.53fF
C255 pd_0/DOWN pd_0/R 0.36fF
C256 pd_0/DIV pd_0/tspc_r_1/z5 0.04fF
C257 pd_0/tspc_r_1/Z1 pd_0/tspc_r_1/Z2 0.71fF
C258 pd_0/tspc_r_1/Z3 pd_0/tspc_r_1/Z4 0.20fF
C259 divider_0/gnd divider_0/nor_1/Z1 0.01fF
C260 ro_complete_0/cbank_0/switch_4/vin ro_complete_0/cbank_0/switch_5/vin 0.19fF
C261 divider_0/prescaler_0/m1_2700_2190# divider_0/prescaler_0/tspc_1/Z3 0.33fF
C262 divider_0/nor_0/Z1 divider_0/nor_0/B 0.06fF
C263 divider_0/vdd divider_0/tspc_2/Z1 0.58fF
C264 divider_0/prescaler_0/Out divider_0/prescaler_0/tspc_1/Z4 0.28fF
C265 ro_complete_0/cbank_2/switch_3/vin ro_complete_0/cbank_2/switch_2/vin 0.20fF
C266 divider_0/tspc_2/Z1 divider_0/tspc_2/Z3 0.06fF
C267 divider_0/nor_1/B divider_0/tspc_2/Z4 0.22fF
C268 pd_0/tspc_r_0/Z3 pd_0/tspc_r_0/Z1 0.09fF
C269 pd_0/REF pd_0/tspc_r_0/Z2 0.19fF
C270 divider_0/mc2 divider_0/prescaler_0/tspc_2/Z2 0.24fF
C271 divider_0/prescaler_0/tspc_0/Z4 divider_0/prescaler_0/tspc_1/Q 0.21fF
C272 divider_0/gnd divider_0/prescaler_0/tspc_2/Q 0.35fF
C273 divider_0/prescaler_0/Out divider_0/vdd 0.75fF
C274 ro_complete_0/a4 ro_complete_0/cbank_1/v 0.05fF
C275 divider_0/tspc_0/Q divider_0/tspc_0/Z3 0.05fF
C276 divider_0/prescaler_0/tspc_2/Z1 divider_0/vdd 0.58fF
C277 divider_0/prescaler_0/tspc_2/Z3 divider_0/prescaler_0/tspc_2/Q 0.05fF
C278 pd_0/tspc_r_0/Qbar pd_0/R 0.03fF
C279 GND pd_0/tspc_r_1/Z2 0.14fF
C280 io_clamp_high[2] io_analog[6] 0.53fF
C281 divider_0/prescaler_0/tspc_0/Z3 divider_0/prescaler_0/tspc_0/Z2 0.16fF
C282 divider_0/prescaler_0/tspc_0/D divider_0/prescaler_0/tspc_1/Q 0.32fF
C283 divider_0/nor_0/A divider_0/vdd 0.83fF
C284 divider_0/vdd divider_0/prescaler_0/tspc_2/D 1.18fF
C285 divider_0/prescaler_0/tspc_2/a_740_n680# divider_0/clk 0.01fF
C286 pd_0/R pd_0/and_pd_0/Out1 0.23fF
C287 ro_complete_0/a3 ro_complete_0/cbank_1/switch_4/vin 0.13fF
C288 ro_complete_0/cbank_0/switch_5/vin ro_complete_0/cbank_0/v 1.30fF
C289 ro_complete_0/cbank_0/switch_2/vin ro_complete_0/a2 0.09fF
C290 divider_0/tspc_1/Z2 divider_0/nor_0/B 0.30fF
C291 divider_0/prescaler_0/Out divider_0/gnd 0.46fF
C292 ro_complete_0/cbank_2/switch_1/vin ro_complete_0/cbank_2/switch_2/vin 0.20fF
C293 divider_0/tspc_0/Z1 divider_0/tspc_0/Z2 1.07fF
C294 divider_0/prescaler_0/tspc_2/Z1 divider_0/prescaler_0/tspc_2/Z3 0.06fF
C295 divider_0/prescaler_0/tspc_2/a_740_n680# divider_0/prescaler_0/tspc_2/a_630_n680# 0.19fF
C296 divider_0/prescaler_0/tspc_1/Z4 divider_0/vdd 0.01fF
C297 divider_0/Out divider_0/tspc_2/a_630_n680# 0.04fF
C298 GND pd_0/tspc_r_0/Z4 0.54fF
C299 divider_0/prescaler_0/tspc_0/Z4 divider_0/prescaler_0/tspc_0/D 0.11fF
C300 divider_0/gnd divider_0/nor_0/A 0.90fF
C301 ro_complete_0/a0 ro_complete_0/cbank_1/switch_1/vin 0.13fF
C302 divider_0/gnd divider_0/prescaler_0/tspc_2/D 0.05fF
C303 divider_0/and_0/A divider_0/and_0/B 0.18fF
C304 divider_0/tspc_1/Z3 divider_0/tspc_1/a_630_n680# 0.05fF
C305 divider_0/prescaler_0/tspc_2/Z3 divider_0/prescaler_0/tspc_2/D 0.05fF
C306 divider_0/prescaler_0/tspc_1/Z2 divider_0/clk 0.11fF
C307 pd_0/tspc_r_1/Qbar1 pd_0/tspc_r_1/z5 0.20fF
C308 divider_0/prescaler_0/tspc_0/Z2 divider_0/prescaler_0/tspc_1/Q 0.06fF
C309 divider_0/prescaler_0/tspc_0/Z1 divider_0/vdd 0.58fF
C310 ro_complete_0/cbank_2/v ro_complete_0/cbank_2/switch_0/vin 1.30fF
C311 divider_0/vdd divider_0/tspc_2/Z3 0.67fF
C312 divider_0/prescaler_0/tspc_2/D divider_0/prescaler_0/nand_1/z1 0.24fF
C313 divider_0/gnd divider_0/prescaler_0/tspc_1/Z4 0.44fF
C314 ro_complete_0/a0 ro_complete_0/cbank_2/v 0.05fF
C315 divider_0/prescaler_0/m1_2700_2190# divider_0/prescaler_0/tspc_1/Q 0.38fF
C316 divider_0/tspc_2/Z1 divider_0/tspc_2/Z4 0.00fF
C317 divider_0/prescaler_0/Out divider_0/tspc_0/Z3 0.45fF
C318 divider_0/gnd divider_0/vdd 0.26fF
C319 ro_complete_0/cbank_0/v ro_complete_0/cbank_2/v 1.27fF
C320 divider_0/tspc_0/a_630_n680# divider_0/tspc_0/Z4 0.12fF
C321 divider_0/prescaler_0/tspc_2/Z3 divider_0/vdd 0.67fF
C322 divider_0/prescaler_0/tspc_0/a_630_n680# divider_0/clk 0.01fF
C323 pd_0/DIV pd_0/tspc_r_1/Qbar1 0.12fF
C324 GND pd_0/R 0.46fF
C325 io_clamp_low[1] io_analog[5] 0.53fF
C326 divider_0/prescaler_0/tspc_0/Z4 divider_0/prescaler_0/tspc_0/Z2 0.36fF
C327 divider_0/gnd divider_0/tspc_2/Z3 0.27fF
C328 divider_0/nor_0/A divider_0/tspc_0/Z3 0.38fF
C329 divider_0/nor_0/B divider_0/tspc_1/Z4 0.21fF
C330 divider_0/vdd divider_0/prescaler_0/nand_1/z1 0.01fF
C331 divider_0/prescaler_0/tspc_0/D divider_0/prescaler_0/tspc_0/Z2 0.09fF
C332 divider_0/tspc_1/Z2 divider_0/tspc_1/Z1 1.07fF
C333 divider_0/tspc_1/Z3 divider_0/tspc_0/Q 0.45fF
C334 divider_0/prescaler_0/tspc_1/Z4 divider_0/prescaler_0/tspc_1/a_630_n680# 0.12fF
C335 divider_0/gnd divider_0/prescaler_0/tspc_2/Z3 0.27fF
C336 ro_complete_0/a2 ro_complete_0/cbank_2/switch_2/vin 0.09fF
C337 divider_0/prescaler_0/tspc_2/Z1 divider_0/prescaler_0/tspc_2/Z4 0.00fF
C338 pd_0/UP pd_0/DOWN 0.46fF
C339 pd_0/tspc_r_0/Z4 pd_0/tspc_r_0/z5 0.04fF
C340 ro_complete_0/cbank_0/switch_1/vin ro_complete_0/cbank_0/switch_2/vin 0.20fF
C341 divider_0/gnd divider_0/prescaler_0/nand_1/z1 0.16fF
C342 ro_complete_0/cbank_2/switch_1/vin ro_complete_0/cbank_2/switch_0/vin 0.20fF
C343 ro_complete_0/cbank_2/switch_4/vin ro_complete_0/cbank_2/v 1.30fF
C344 divider_0/vdd divider_0/tspc_0/Z3 0.67fF
C345 divider_0/prescaler_0/tspc_1/Q divider_0/prescaler_0/nand_0/z1 0.22fF
C346 divider_0/prescaler_0/tspc_2/Z4 divider_0/prescaler_0/tspc_2/D 0.11fF
C347 ro_complete_0/cbank_0/switch_1/vin ro_complete_0/cbank_0/switch_0/vin 0.20fF
C348 divider_0/prescaler_0/tspc_1/Z1 divider_0/prescaler_0/tspc_1/Z2 1.07fF
C349 divider_0/nor_0/B divider_0/and_0/B 0.35fF
C350 divider_0/vdd divider_0/tspc_2/Z4 0.01fF
C351 divider_0/prescaler_0/tspc_2/Q divider_0/clk 0.05fF
C352 divider_0/gnd divider_0/prescaler_0/tspc_1/a_630_n680# 0.61fF
C353 ro_complete_0/a3 ro_complete_0/cbank_1/v 0.05fF
C354 ro_complete_0/cbank_2/switch_3/vin ro_complete_0/cbank_2/switch_4/vin 0.20fF
C355 divider_0/tspc_0/a_630_n680# divider_0/tspc_0/Q 0.04fF
C356 divider_0/and_0/OUT divider_0/and_0/B 0.01fF
C357 divider_0/tspc_2/Z3 divider_0/tspc_2/Z4 0.65fF
C358 pd_0/tspc_r_0/Z3 GND 0.32fF
C359 pd_0/REF pd_0/tspc_r_0/Z4 0.02fF
C360 pd_0/UP pd_0/tspc_r_0/Qbar 0.21fF
C361 divider_0/gnd divider_0/tspc_0/Z3 0.27fF
C362 divider_0/prescaler_0/tspc_2/Z4 divider_0/vdd 0.01fF
C363 divider_0/prescaler_0/tspc_2/a_630_n680# divider_0/prescaler_0/tspc_2/Q 0.04fF
C364 pd_0/UP pd_0/and_pd_0/Out1 0.13fF
C365 pd_0/tspc_r_1/Z3 pd_0/DOWN 0.03fF
C366 GND pd_0/tspc_r_1/Z4 0.54fF
C367 ro_complete_0/cbank_0/switch_3/vin ro_complete_0/a3 0.09fF
C368 divider_0/gnd divider_0/tspc_2/Z4 0.44fF
C369 divider_0/prescaler_0/tspc_0/D divider_0/prescaler_0/nand_0/z1 0.21fF
C370 divider_0/prescaler_0/Out divider_0/clk 0.51fF
C371 divider_0/tspc_1/Z1 divider_0/tspc_1/Z4 0.00fF
C372 divider_0/nor_0/B divider_0/tspc_1/a_630_n680# 0.35fF
C373 pd_0/R pd_0/and_pd_0/Z1 0.02fF
C374 divider_0/vdd divider_0/and_0/out1 1.44fF
C375 divider_0/prescaler_0/tspc_2/D divider_0/clk 0.26fF
C376 divider_0/gnd divider_0/prescaler_0/tspc_2/Z4 0.44fF
C377 ro_complete_0/a1 ro_complete_0/cbank_1/v 0.05fF
C378 divider_0/prescaler_0/tspc_1/Z2 divider_0/and_0/OUT 0.06fF
C379 divider_0/prescaler_0/tspc_2/Z3 divider_0/prescaler_0/tspc_2/Z4 0.65fF
C380 cp_0/a_1710_n2840# cp_0/out 0.61fF
C381 pd_0/REF pd_0/R 0.61fF
C382 divider_0/nor_0/B divider_0/nor_1/B 0.48fF
C383 divider_0/prescaler_0/tspc_1/Z4 divider_0/clk 0.12fF
C384 divider_0/and_0/B divider_0/and_0/Z1 0.07fF
C385 divider_0/gnd divider_0/and_0/out1 0.23fF
C386 divider_0/prescaler_0/tspc_1/Z2 divider_0/prescaler_0/tspc_1/Z3 0.16fF
C387 divider_0/vdd divider_0/clk 0.27fF
C388 divider_0/prescaler_0/Out divider_0/tspc_0/a_630_n680# 0.01fF
C389 divider_0/nor_0/A divider_0/and_0/A 0.01fF
C390 ro_complete_0/cbank_0/switch_5/vin ro_complete_0/a5 0.09fF
C391 divider_0/tspc_1/Z3 divider_0/vdd 0.67fF
C392 divider_0/nor_0/B divider_0/tspc_0/Q 0.22fF
C393 divider_0/tspc_1/Q divider_0/tspc_1/a_630_n680# 0.04fF
C394 pd_0/tspc_r_0/Z3 pd_0/tspc_r_0/z5 0.11fF
C395 pd_0/UP GND 0.26fF
C396 divider_0/nor_0/A divider_0/tspc_0/a_630_n680# 0.35fF
C397 pd_0/tspc_r_1/Z3 pd_0/tspc_r_1/Z1 0.09fF
C398 pd_0/DIV pd_0/tspc_r_1/Z2 0.19fF
C399 io_clamp_high[0] io_analog[4] 0.53fF
C400 divider_0/nor_1/Z1 divider_0/nor_0/B 0.26fF
C401 divider_0/gnd divider_0/clk 0.07fF
C402 divider_0/prescaler_0/tspc_2/Z3 divider_0/clk 0.45fF
C403 divider_0/gnd divider_0/tspc_1/Z3 0.27fF
C404 divider_0/prescaler_0/Out divider_0/prescaler_0/tspc_1/Z1 0.08fF
C405 ro_complete_0/a0 ro_complete_0/cbank_1/switch_0/vin 0.09fF
C406 divider_0/mc2 divider_0/and_0/B 0.20fF
C407 divider_0/and_0/A divider_0/vdd 0.11fF
C408 divider_0/nor_1/B divider_0/tspc_1/Q 0.22fF
C409 pd_0/REF pd_0/tspc_r_0/Z3 0.65fF
C410 divider_0/prescaler_0/tspc_0/a_740_n680# divider_0/prescaler_0/tspc_1/Z2 0.01fF
C411 divider_0/gnd divider_0/prescaler_0/tspc_2/a_630_n680# 0.61fF
C412 ro_complete_0/cbank_2/switch_3/vin ro_complete_0/cbank_2/v 1.30fF
C413 ro_complete_0/cbank_1/switch_5/vin ro_complete_0/a5 0.09fF
C414 divider_0/tspc_0/Z1 divider_0/tspc_0/Z4 0.00fF
C415 divider_0/prescaler_0/tspc_2/Z3 divider_0/prescaler_0/tspc_2/a_630_n680# 0.05fF
C416 cp_0/upbar cp_0/down 0.02fF
C417 pd_0/tspc_r_0/Qbar pd_0/DOWN 0.02fF
C418 GND pd_0/tspc_r_1/Z3 0.32fF
C419 pd_0/tspc_r_0/Qbar1 pd_0/R 0.30fF
C420 ro_complete_0/cbank_0/switch_3/vin ro_complete_0/cbank_0/switch_2/vin 0.20fF
C421 ro_complete_0/a5 ro_complete_0/cbank_2/v 0.10fF
C422 divider_0/prescaler_0/tspc_2/Q divider_0/and_0/OUT 0.04fF
C423 divider_0/prescaler_0/tspc_1/a_630_n680# divider_0/clk 0.01fF
C424 divider_0/prescaler_0/tspc_0/Z3 divider_0/prescaler_0/tspc_0/a_630_n680# 0.05fF
C425 divider_0/gnd divider_0/and_0/A 0.53fF
C426 divider_0/prescaler_0/tspc_1/Z1 divider_0/prescaler_0/tspc_1/Z4 0.00fF
C427 divider_0/gnd divider_0/tspc_0/a_630_n680# 0.62fF
C428 divider_0/prescaler_0/tspc_0/a_740_n680# divider_0/prescaler_0/tspc_0/a_630_n680# 0.19fF
C429 divider_0/tspc_0/Q divider_0/tspc_1/Z1 0.01fF
C430 divider_0/prescaler_0/tspc_1/Z2 divider_0/prescaler_0/tspc_1/Q 0.06fF
C431 divider_0/prescaler_0/tspc_1/Z1 divider_0/vdd 0.58fF
C432 divider_0/nor_1/B divider_0/tspc_2/a_630_n680# 0.35fF
C433 pd_0/UP pd_0/tspc_r_0/z5 0.03fF
C434 ro_complete_0/cbank_0/switch_1/vin ro_complete_0/a0 0.13fF
C435 divider_0/nor_0/A divider_0/nor_0/B 1.22fF
C436 ro_complete_0/cbank_2/switch_1/vin ro_complete_0/cbank_2/v 1.30fF
C437 pd_0/tspc_r_0/Qbar pd_0/and_pd_0/Out1 0.05fF
C438 pd_0/UP pd_0/and_pd_0/Z1 0.06fF
C439 pd_0/DIV pd_0/R 0.51fF
C440 ro_complete_0/cbank_1/switch_1/vin ro_complete_0/cbank_1/switch_2/vin 0.20fF
C441 ro_complete_0/cbank_0/switch_1/vin ro_complete_0/cbank_0/v 1.30fF
C442 divider_0/mc2 divider_0/nor_1/B 0.15fF
C443 divider_0/and_0/OUT divider_0/prescaler_0/tspc_2/D 0.03fF
C444 divider_0/prescaler_0/tspc_2/Z4 divider_0/clk 0.12fF
C445 divider_0/prescaler_0/Out divider_0/prescaler_0/tspc_1/Z3 0.11fF
C446 ro_complete_0/cbank_0/switch_4/vin ro_complete_0/a4 0.09fF
C447 divider_0/tspc_1/Q divider_0/tspc_2/Z1 0.01fF
C448 divider_0/nor_1/B divider_0/tspc_2/Z2 0.40fF
C449 cp_0/a_1710_0# cp_0/a_1710_n2840# 0.83fF
C450 pd_0/tspc_r_0/Z3 pd_0/tspc_r_0/Qbar1 0.38fF
C451 divider_0/nor_0/B divider_0/vdd 0.30fF
C452 divider_0/tspc_0/a_630_n680# divider_0/tspc_0/Z3 0.05fF
C453 divider_0/prescaler_0/tspc_2/Z4 divider_0/prescaler_0/tspc_2/a_630_n680# 0.12fF
C454 GND pd_0/DOWN 0.79fF
C455 divider_0/tspc_0/Z2 divider_0/tspc_0/Z4 0.36fF
C456 divider_0/vdd divider_0/and_0/OUT 1.59fF
C457 pd_0/tspc_r_1/Z4 pd_0/tspc_r_1/z5 0.04fF
C458 divider_0/prescaler_0/tspc_0/Z4 divider_0/prescaler_0/tspc_0/a_630_n680# 0.12fF
C459 ro_complete_0/cbank_0/switch_2/vin ro_complete_0/a1 0.14fF
C460 divider_0/prescaler_0/tspc_1/Z3 divider_0/prescaler_0/tspc_1/Z4 0.65fF
C461 divider_0/prescaler_0/tspc_0/Z3 divider_0/prescaler_0/Out 0.05fF
C462 divider_0/gnd divider_0/nor_0/B 0.99fF
C463 divider_0/prescaler_0/tspc_1/Z3 divider_0/vdd 0.67fF
C464 pd_0/tspc_r_0/Qbar GND 0.18fF
C465 pd_0/tspc_r_0/Z2 pd_0/tspc_r_0/Z4 0.14fF
C466 divider_0/prescaler_0/Out divider_0/prescaler_0/tspc_0/a_740_n680# 0.21fF
C467 divider_0/gnd divider_0/and_0/OUT 0.26fF
C468 ro_complete_0/a2 ro_complete_0/cbank_2/v 0.05fF
C469 divider_0/nor_0/Z1 divider_0/and_0/B 0.18fF
C470 divider_0/and_0/A divider_0/and_0/out1 0.01fF
C471 divider_0/tspc_1/Z2 divider_0/tspc_1/Z4 0.36fF
C472 divider_0/prescaler_0/tspc_2/Q divider_0/prescaler_0/tspc_1/Q 0.19fF
C473 GND pd_0/and_pd_0/Out1 0.18fF
C474 pd_0/tspc_r_1/Qbar1 pd_0/R 0.01fF
C475 pd_0/DIV pd_0/tspc_r_1/Z4 0.02fF
C476 pd_0/DOWN pd_0/tspc_r_1/Qbar 0.21fF
C477 divider_0/vdd divider_0/tspc_1/Q 0.72fF
C478 divider_0/and_0/OUT divider_0/prescaler_0/nand_1/z1 0.01fF
C479 divider_0/prescaler_0/tspc_2/a_630_n680# divider_0/clk 0.01fF
C480 divider_0/gnd divider_0/prescaler_0/tspc_1/Z3 0.27fF
C481 ro_complete_0/cbank_1/switch_1/vin ro_complete_0/cbank_1/switch_0/vin 0.20fF
C482 io_analog[4] vdd 25.05fF
C483 io_analog[5] vdd 25.05fF
C484 io_analog[6] vdd 25.05fF
C485 io_in_3v3[0] vdd 0.61fF
C486 io_oeb[26] vdd 0.61fF
C487 io_in[0] vdd 0.61fF
C488 io_out[26] vdd 0.61fF
C489 io_out[0] vdd 0.61fF
C490 io_in[26] vdd 0.61fF
C491 io_oeb[0] vdd 0.61fF
C492 io_in_3v3[26] vdd 0.61fF
C493 io_in_3v3[1] vdd 0.61fF
C494 io_oeb[25] vdd 0.61fF
C495 io_in[1] vdd 0.61fF
C496 io_out[25] vdd 0.61fF
C497 io_out[1] vdd 0.61fF
C498 io_in[25] vdd 0.61fF
C499 io_oeb[1] vdd 0.61fF
C500 io_in_3v3[25] vdd 0.61fF
C501 io_in_3v3[2] vdd 0.61fF
C502 io_oeb[24] vdd 0.61fF
C503 io_in[2] vdd 0.61fF
C504 io_out[24] vdd 0.61fF
C505 io_out[2] vdd 0.61fF
C506 io_in[24] vdd 0.61fF
C507 io_oeb[2] vdd 0.61fF
C508 io_in_3v3[24] vdd 0.61fF
C509 io_in_3v3[3] vdd 0.61fF
C510 gpio_noesd[17] vdd 0.61fF
C511 io_in[3] vdd 0.61fF
C512 gpio_analog[17] vdd 0.61fF
C513 io_out[3] vdd 0.61fF
C514 io_oeb[3] vdd 0.61fF
C515 io_in_3v3[4] vdd 0.61fF
C516 io_in[4] vdd 0.61fF
C517 io_out[4] vdd 0.61fF
C518 io_oeb[4] vdd 0.61fF
C519 io_oeb[23] vdd 0.61fF
C520 io_out[23] vdd 0.61fF
C521 io_in[23] vdd 0.61fF
C522 io_in_3v3[23] vdd 0.61fF
C523 gpio_noesd[16] vdd 0.61fF
C524 gpio_analog[16] vdd 0.61fF
C525 io_in_3v3[5] vdd 0.61fF
C526 io_in[5] vdd 0.61fF
C527 io_out[5] vdd 0.61fF
C528 io_oeb[5] vdd 0.61fF
C529 io_oeb[22] vdd 0.61fF
C530 io_out[22] vdd 0.61fF
C531 io_in[22] vdd 0.61fF
C532 io_in_3v3[22] vdd 0.61fF
C533 gpio_noesd[15] vdd 0.61fF
C534 gpio_analog[15] vdd 0.61fF
C535 io_in_3v3[6] vdd 0.61fF
C536 io_in[6] vdd 0.61fF
C537 io_out[6] vdd 0.61fF
C538 io_oeb[6] vdd 0.61fF
C539 io_oeb[21] vdd 0.61fF
C540 io_out[21] vdd 0.61fF
C541 io_in[21] vdd 0.61fF
C542 io_in_3v3[21] vdd 0.61fF
C543 gpio_noesd[14] vdd 0.61fF
C544 gpio_analog[14] vdd 0.61fF
C545 vssa1 vdd 26.08fF
C546 vssd2 vdd 13.04fF
C547 vssd1 vdd 13.04fF
C548 vdda2 vdd 13.04fF
C549 vdda1 vdd 26.08fF
C550 io_oeb[20] vdd 0.61fF
C551 io_out[20] vdd 0.61fF
C552 io_in[20] vdd 0.61fF
C553 io_in_3v3[20] vdd 0.61fF
C554 gpio_noesd[13] vdd 0.61fF
C555 gpio_analog[13] vdd 0.61fF
C556 gpio_analog[0] vdd 0.61fF
C557 gpio_noesd[0] vdd 0.61fF
C558 io_in_3v3[7] vdd 0.61fF
C559 io_in[7] vdd 0.61fF
C560 io_out[7] vdd 0.61fF
C561 io_oeb[7] vdd 0.61fF
C562 io_oeb[19] vdd 0.61fF
C563 io_out[19] vdd 0.61fF
C564 io_in[19] vdd 0.61fF
C565 io_in_3v3[19] vdd 0.61fF
C566 gpio_noesd[12] vdd 0.61fF
C567 gpio_analog[12] vdd 0.61fF
C568 gpio_analog[1] vdd 0.61fF
C569 gpio_noesd[1] vdd 0.61fF
C570 io_in_3v3[8] vdd 0.61fF
C571 io_in[8] vdd 0.61fF
C572 io_out[8] vdd 0.61fF
C573 io_oeb[8] vdd 0.61fF
C574 io_oeb[18] vdd 0.61fF
C575 io_out[18] vdd 0.61fF
C576 io_in[18] vdd 0.61fF
C577 io_in_3v3[18] vdd 0.61fF
C578 gpio_noesd[11] vdd 0.61fF
C579 gpio_analog[11] vdd 0.61fF
C580 gpio_analog[2] vdd 0.61fF
C581 gpio_noesd[2] vdd 0.61fF
C582 io_in_3v3[9] vdd 0.61fF
C583 io_in[9] vdd 0.61fF
C584 io_out[9] vdd 0.61fF
C585 io_oeb[9] vdd 0.61fF
C586 io_oeb[17] vdd 0.61fF
C587 io_out[17] vdd 0.61fF
C588 io_in[17] vdd 0.61fF
C589 io_in_3v3[17] vdd 0.61fF
C590 gpio_noesd[10] vdd 0.61fF
C591 gpio_analog[10] vdd 0.61fF
C592 gpio_analog[3] vdd 0.61fF
C593 gpio_noesd[3] vdd 0.61fF
C594 io_in_3v3[10] vdd 0.61fF
C595 io_in[10] vdd 0.61fF
C596 io_out[10] vdd 0.61fF
C597 io_oeb[10] vdd 0.61fF
C598 io_oeb[16] vdd 0.61fF
C599 io_out[16] vdd 0.61fF
C600 io_in[16] vdd 0.61fF
C601 io_in_3v3[16] vdd 0.61fF
C602 gpio_noesd[9] vdd 0.61fF
C603 gpio_analog[9] vdd 0.61fF
C604 gpio_analog[4] vdd 0.61fF
C605 gpio_noesd[4] vdd 0.61fF
C606 io_in_3v3[11] vdd 0.61fF
C607 io_in[11] vdd 0.61fF
C608 io_out[11] vdd 0.61fF
C609 io_oeb[11] vdd 0.61fF
C610 io_oeb[15] vdd 0.61fF
C611 io_out[15] vdd 0.61fF
C612 io_in[15] vdd 0.61fF
C613 io_in_3v3[15] vdd 0.61fF
C614 gpio_noesd[8] vdd 0.61fF
C615 gpio_analog[8] vdd 0.61fF
C616 gpio_analog[5] vdd 0.61fF
C617 gpio_noesd[5] vdd 0.61fF
C618 io_in_3v3[12] vdd 0.61fF
C619 io_in[12] vdd 0.61fF
C620 io_out[12] vdd 0.61fF
C621 io_oeb[12] vdd 0.61fF
C622 io_oeb[14] vdd 0.61fF
C623 io_out[14] vdd 0.61fF
C624 io_in[14] vdd 0.61fF
C625 io_in_3v3[14] vdd 0.61fF
C626 gpio_noesd[7] vdd 0.61fF
C627 gpio_analog[7] vdd 0.61fF
C628 vssa2 vdd 13.04fF
C629 gpio_analog[6] vdd 0.61fF
C630 gpio_noesd[6] vdd 0.61fF
C631 io_in_3v3[13] vdd 0.61fF
C632 io_in[13] vdd 0.61fF
C633 io_out[13] vdd 0.61fF
C634 io_oeb[13] vdd 0.61fF
C635 vccd1 vdd 13.04fF
C636 vccd2 vdd 13.04fF
C637 io_analog[0] vdd 6.83fF
C638 io_analog[10] vdd 6.83fF
C639 io_analog[1] vdd 6.83fF
C640 io_analog[2] vdd 6.83fF
C641 io_analog[3] vdd 6.83fF
C642 io_clamp_high[0] vdd 3.58fF
C643 io_clamp_low[0] vdd 3.58fF
C644 io_clamp_high[1] vdd 3.58fF
C645 io_clamp_low[1] vdd 3.58fF
C646 io_clamp_high[2] vdd 3.58fF
C647 io_clamp_low[2] vdd 3.58fF
C648 io_analog[7] vdd 6.83fF
C649 io_analog[8] vdd 6.83fF
C650 io_analog[9] vdd 6.83fF
C651 user_irq[2] vdd 0.63fF
C652 user_irq[1] vdd 0.63fF
C653 user_irq[0] vdd 0.63fF
C654 user_clock2 vdd 0.63fF
C655 la_oenb[127] vdd 0.63fF
C656 la_data_out[127] vdd 0.63fF
C657 la_data_in[127] vdd 0.63fF
C658 la_oenb[126] vdd 0.63fF
C659 la_data_out[126] vdd 0.63fF
C660 la_data_in[126] vdd 0.63fF
C661 la_oenb[125] vdd 0.63fF
C662 la_data_out[125] vdd 0.63fF
C663 la_data_in[125] vdd 0.63fF
C664 la_oenb[124] vdd 0.63fF
C665 la_data_out[124] vdd 0.63fF
C666 la_data_in[124] vdd 0.63fF
C667 la_oenb[123] vdd 0.63fF
C668 la_data_out[123] vdd 0.63fF
C669 la_data_in[123] vdd 0.63fF
C670 la_oenb[122] vdd 0.63fF
C671 la_data_out[122] vdd 0.63fF
C672 la_data_in[122] vdd 0.63fF
C673 la_oenb[121] vdd 0.63fF
C674 la_data_out[121] vdd 0.63fF
C675 la_data_in[121] vdd 0.63fF
C676 la_oenb[120] vdd 0.63fF
C677 la_data_out[120] vdd 0.63fF
C678 la_data_in[120] vdd 0.63fF
C679 la_oenb[119] vdd 0.63fF
C680 la_data_out[119] vdd 0.63fF
C681 la_data_in[119] vdd 0.63fF
C682 la_oenb[118] vdd 0.63fF
C683 la_data_out[118] vdd 0.63fF
C684 la_data_in[118] vdd 0.63fF
C685 la_oenb[117] vdd 0.63fF
C686 la_data_out[117] vdd 0.63fF
C687 la_data_in[117] vdd 0.63fF
C688 la_oenb[116] vdd 0.63fF
C689 la_data_out[116] vdd 0.63fF
C690 la_data_in[116] vdd 0.63fF
C691 la_oenb[115] vdd 0.63fF
C692 la_data_out[115] vdd 0.63fF
C693 la_data_in[115] vdd 0.63fF
C694 la_oenb[114] vdd 0.63fF
C695 la_data_out[114] vdd 0.63fF
C696 la_data_in[114] vdd 0.63fF
C697 la_oenb[113] vdd 0.63fF
C698 la_data_out[113] vdd 0.63fF
C699 la_data_in[113] vdd 0.63fF
C700 la_oenb[112] vdd 0.63fF
C701 la_data_out[112] vdd 0.63fF
C702 la_data_in[112] vdd 0.63fF
C703 la_oenb[111] vdd 0.63fF
C704 la_data_out[111] vdd 0.63fF
C705 la_data_in[111] vdd 0.63fF
C706 la_oenb[110] vdd 0.63fF
C707 la_data_out[110] vdd 0.63fF
C708 la_data_in[110] vdd 0.63fF
C709 la_oenb[109] vdd 0.63fF
C710 la_data_out[109] vdd 0.63fF
C711 la_data_in[109] vdd 0.63fF
C712 la_oenb[108] vdd 0.63fF
C713 la_data_out[108] vdd 0.63fF
C714 la_data_in[108] vdd 0.63fF
C715 la_oenb[107] vdd 0.63fF
C716 la_data_out[107] vdd 0.63fF
C717 la_data_in[107] vdd 0.63fF
C718 la_oenb[106] vdd 0.63fF
C719 la_data_out[106] vdd 0.63fF
C720 la_data_in[106] vdd 0.63fF
C721 la_oenb[105] vdd 0.63fF
C722 la_data_out[105] vdd 0.63fF
C723 la_data_in[105] vdd 0.63fF
C724 la_oenb[104] vdd 0.63fF
C725 la_data_out[104] vdd 0.63fF
C726 la_data_in[104] vdd 0.63fF
C727 la_oenb[103] vdd 0.63fF
C728 la_data_out[103] vdd 0.63fF
C729 la_data_in[103] vdd 0.63fF
C730 la_oenb[102] vdd 0.63fF
C731 la_data_out[102] vdd 0.63fF
C732 la_data_in[102] vdd 0.63fF
C733 la_oenb[101] vdd 0.63fF
C734 la_data_out[101] vdd 0.63fF
C735 la_data_in[101] vdd 0.63fF
C736 la_oenb[100] vdd 0.63fF
C737 la_data_out[100] vdd 0.63fF
C738 la_data_in[100] vdd 0.63fF
C739 la_oenb[99] vdd 0.63fF
C740 la_data_out[99] vdd 0.63fF
C741 la_data_in[99] vdd 0.63fF
C742 la_oenb[98] vdd 0.63fF
C743 la_data_out[98] vdd 0.63fF
C744 la_data_in[98] vdd 0.63fF
C745 la_oenb[97] vdd 0.63fF
C746 la_data_out[97] vdd 0.63fF
C747 la_data_in[97] vdd 0.63fF
C748 la_oenb[96] vdd 0.63fF
C749 la_data_out[96] vdd 0.63fF
C750 la_data_in[96] vdd 0.63fF
C751 la_oenb[95] vdd 0.63fF
C752 la_data_out[95] vdd 0.63fF
C753 la_data_in[95] vdd 0.63fF
C754 la_oenb[94] vdd 0.63fF
C755 la_data_out[94] vdd 0.63fF
C756 la_data_in[94] vdd 0.63fF
C757 la_oenb[93] vdd 0.63fF
C758 la_data_out[93] vdd 0.63fF
C759 la_data_in[93] vdd 0.63fF
C760 la_oenb[92] vdd 0.63fF
C761 la_data_out[92] vdd 0.63fF
C762 la_data_in[92] vdd 0.63fF
C763 la_oenb[91] vdd 0.63fF
C764 la_data_out[91] vdd 0.63fF
C765 la_data_in[91] vdd 0.63fF
C766 la_oenb[90] vdd 0.63fF
C767 la_data_out[90] vdd 0.63fF
C768 la_data_in[90] vdd 0.63fF
C769 la_oenb[89] vdd 0.63fF
C770 la_data_out[89] vdd 0.63fF
C771 la_data_in[89] vdd 0.63fF
C772 la_oenb[88] vdd 0.63fF
C773 la_data_out[88] vdd 0.63fF
C774 la_data_in[88] vdd 0.63fF
C775 la_oenb[87] vdd 0.63fF
C776 la_data_out[87] vdd 0.63fF
C777 la_data_in[87] vdd 0.63fF
C778 la_oenb[86] vdd 0.63fF
C779 la_data_out[86] vdd 0.63fF
C780 la_data_in[86] vdd 0.63fF
C781 la_oenb[85] vdd 0.63fF
C782 la_data_out[85] vdd 0.63fF
C783 la_data_in[85] vdd 0.63fF
C784 la_oenb[84] vdd 0.63fF
C785 la_data_out[84] vdd 0.63fF
C786 la_data_in[84] vdd 0.63fF
C787 la_oenb[83] vdd 0.63fF
C788 la_data_out[83] vdd 0.63fF
C789 la_data_in[83] vdd 0.63fF
C790 la_oenb[82] vdd 0.63fF
C791 la_data_out[82] vdd 0.63fF
C792 la_data_in[82] vdd 0.63fF
C793 la_oenb[81] vdd 0.63fF
C794 la_data_out[81] vdd 0.63fF
C795 la_data_in[81] vdd 0.63fF
C796 la_oenb[80] vdd 0.63fF
C797 la_data_out[80] vdd 0.63fF
C798 la_data_in[80] vdd 0.63fF
C799 la_oenb[79] vdd 0.63fF
C800 la_data_out[79] vdd 0.63fF
C801 la_data_in[79] vdd 0.63fF
C802 la_oenb[78] vdd 0.63fF
C803 la_data_out[78] vdd 0.63fF
C804 la_data_in[78] vdd 0.63fF
C805 la_oenb[77] vdd 0.63fF
C806 la_data_out[77] vdd 0.63fF
C807 la_data_in[77] vdd 0.63fF
C808 la_oenb[76] vdd 0.63fF
C809 la_data_out[76] vdd 0.63fF
C810 la_data_in[76] vdd 0.63fF
C811 la_oenb[75] vdd 0.63fF
C812 la_data_out[75] vdd 0.63fF
C813 la_data_in[75] vdd 0.63fF
C814 la_oenb[74] vdd 0.63fF
C815 la_data_out[74] vdd 0.63fF
C816 la_data_in[74] vdd 0.63fF
C817 la_oenb[73] vdd 0.63fF
C818 la_data_out[73] vdd 0.63fF
C819 la_data_in[73] vdd 0.63fF
C820 la_oenb[72] vdd 0.63fF
C821 la_data_out[72] vdd 0.63fF
C822 la_data_in[72] vdd 0.63fF
C823 la_oenb[71] vdd 0.63fF
C824 la_data_out[71] vdd 0.63fF
C825 la_data_in[71] vdd 0.63fF
C826 la_oenb[70] vdd 0.63fF
C827 la_data_out[70] vdd 0.63fF
C828 la_data_in[70] vdd 0.63fF
C829 la_oenb[69] vdd 0.63fF
C830 la_data_out[69] vdd 0.63fF
C831 la_data_in[69] vdd 0.63fF
C832 la_oenb[68] vdd 0.63fF
C833 la_data_out[68] vdd 0.63fF
C834 la_data_in[68] vdd 0.63fF
C835 la_oenb[67] vdd 0.63fF
C836 la_data_out[67] vdd 0.63fF
C837 la_data_in[67] vdd 0.63fF
C838 la_oenb[66] vdd 0.63fF
C839 la_data_out[66] vdd 0.63fF
C840 la_data_in[66] vdd 0.63fF
C841 la_oenb[65] vdd 0.63fF
C842 la_data_out[65] vdd 0.63fF
C843 la_data_in[65] vdd 0.63fF
C844 la_oenb[64] vdd 0.63fF
C845 la_data_out[64] vdd 0.63fF
C846 la_data_in[64] vdd 0.63fF
C847 la_oenb[63] vdd 0.63fF
C848 la_data_out[63] vdd 0.63fF
C849 la_data_in[63] vdd 0.63fF
C850 la_oenb[62] vdd 0.63fF
C851 la_data_out[62] vdd 0.63fF
C852 la_data_in[62] vdd 0.63fF
C853 la_oenb[61] vdd 0.63fF
C854 la_data_out[61] vdd 0.63fF
C855 la_data_in[61] vdd 0.63fF
C856 la_oenb[60] vdd 0.63fF
C857 la_data_out[60] vdd 0.63fF
C858 la_data_in[60] vdd 0.63fF
C859 la_oenb[59] vdd 0.63fF
C860 la_data_out[59] vdd 0.63fF
C861 la_data_in[59] vdd 0.63fF
C862 la_oenb[58] vdd 0.63fF
C863 la_data_out[58] vdd 0.63fF
C864 la_data_in[58] vdd 0.63fF
C865 la_oenb[57] vdd 0.63fF
C866 la_data_out[57] vdd 0.63fF
C867 la_data_in[57] vdd 0.63fF
C868 la_oenb[56] vdd 0.63fF
C869 la_data_out[56] vdd 0.63fF
C870 la_data_in[56] vdd 0.63fF
C871 la_oenb[55] vdd 0.63fF
C872 la_data_out[55] vdd 0.63fF
C873 la_data_in[55] vdd 0.63fF
C874 la_oenb[54] vdd 0.63fF
C875 la_data_out[54] vdd 0.63fF
C876 la_data_in[54] vdd 0.63fF
C877 la_oenb[53] vdd 0.63fF
C878 la_data_out[53] vdd 0.63fF
C879 la_data_in[53] vdd 0.63fF
C880 la_oenb[52] vdd 0.63fF
C881 la_data_out[52] vdd 0.63fF
C882 la_data_in[52] vdd 0.63fF
C883 la_oenb[51] vdd 0.63fF
C884 la_data_out[51] vdd 0.63fF
C885 la_data_in[51] vdd 0.63fF
C886 la_oenb[50] vdd 0.63fF
C887 la_data_out[50] vdd 0.63fF
C888 la_data_in[50] vdd 0.63fF
C889 la_oenb[49] vdd 0.63fF
C890 la_data_out[49] vdd 0.63fF
C891 la_data_in[49] vdd 0.63fF
C892 la_oenb[48] vdd 0.63fF
C893 la_data_out[48] vdd 0.63fF
C894 la_data_in[48] vdd 0.63fF
C895 la_oenb[47] vdd 0.63fF
C896 la_data_out[47] vdd 0.63fF
C897 la_data_in[47] vdd 0.63fF
C898 la_oenb[46] vdd 0.63fF
C899 la_data_out[46] vdd 0.63fF
C900 la_data_in[46] vdd 0.63fF
C901 la_oenb[45] vdd 0.63fF
C902 la_data_out[45] vdd 0.63fF
C903 la_data_in[45] vdd 0.63fF
C904 la_oenb[44] vdd 0.63fF
C905 la_data_out[44] vdd 0.63fF
C906 la_data_in[44] vdd 0.63fF
C907 la_oenb[43] vdd 0.63fF
C908 la_data_out[43] vdd 0.63fF
C909 la_data_in[43] vdd 0.63fF
C910 la_oenb[42] vdd 0.63fF
C911 la_data_out[42] vdd 0.63fF
C912 la_data_in[42] vdd 0.63fF
C913 la_oenb[41] vdd 0.63fF
C914 la_data_out[41] vdd 0.63fF
C915 la_data_in[41] vdd 0.63fF
C916 la_oenb[40] vdd 0.63fF
C917 la_data_out[40] vdd 0.63fF
C918 la_data_in[40] vdd 0.63fF
C919 la_oenb[39] vdd 0.63fF
C920 la_data_out[39] vdd 0.63fF
C921 la_data_in[39] vdd 0.63fF
C922 la_oenb[38] vdd 0.63fF
C923 la_data_out[38] vdd 0.63fF
C924 la_data_in[38] vdd 0.63fF
C925 la_oenb[37] vdd 0.63fF
C926 la_data_out[37] vdd 0.63fF
C927 la_data_in[37] vdd 0.63fF
C928 la_oenb[36] vdd 0.63fF
C929 la_data_out[36] vdd 0.63fF
C930 la_data_in[36] vdd 0.63fF
C931 la_oenb[35] vdd 0.63fF
C932 la_data_out[35] vdd 0.63fF
C933 la_data_in[35] vdd 0.63fF
C934 la_oenb[34] vdd 0.63fF
C935 la_data_out[34] vdd 0.63fF
C936 la_data_in[34] vdd 0.63fF
C937 la_oenb[33] vdd 0.63fF
C938 la_data_out[33] vdd 0.63fF
C939 la_data_in[33] vdd 0.63fF
C940 la_oenb[32] vdd 0.63fF
C941 la_data_out[32] vdd 0.63fF
C942 la_data_in[32] vdd 0.63fF
C943 la_oenb[31] vdd 0.63fF
C944 la_data_out[31] vdd 0.63fF
C945 la_data_in[31] vdd 0.63fF
C946 la_oenb[30] vdd 0.63fF
C947 la_data_out[30] vdd 0.63fF
C948 la_data_in[30] vdd 0.63fF
C949 la_oenb[29] vdd 0.63fF
C950 la_data_out[29] vdd 0.63fF
C951 la_data_in[29] vdd 0.63fF
C952 la_oenb[28] vdd 0.63fF
C953 la_data_out[28] vdd 0.63fF
C954 la_data_in[28] vdd 0.63fF
C955 la_oenb[27] vdd 0.63fF
C956 la_data_out[27] vdd 0.63fF
C957 la_data_in[27] vdd 0.63fF
C958 la_oenb[26] vdd 0.63fF
C959 la_data_out[26] vdd 0.63fF
C960 la_data_in[26] vdd 0.63fF
C961 la_oenb[25] vdd 0.63fF
C962 la_data_out[25] vdd 0.63fF
C963 la_data_in[25] vdd 0.63fF
C964 la_oenb[24] vdd 0.63fF
C965 la_data_out[24] vdd 0.63fF
C966 la_data_in[24] vdd 0.63fF
C967 la_oenb[23] vdd 0.63fF
C968 la_data_out[23] vdd 0.63fF
C969 la_data_in[23] vdd 0.63fF
C970 la_oenb[22] vdd 0.63fF
C971 la_data_out[22] vdd 0.63fF
C972 la_data_in[22] vdd 0.63fF
C973 la_oenb[21] vdd 0.63fF
C974 la_data_out[21] vdd 0.63fF
C975 la_data_in[21] vdd 0.63fF
C976 la_oenb[20] vdd 0.63fF
C977 la_data_out[20] vdd 0.63fF
C978 la_data_in[20] vdd 0.63fF
C979 la_oenb[19] vdd 0.63fF
C980 la_data_out[19] vdd 0.63fF
C981 la_data_in[19] vdd 0.63fF
C982 la_oenb[18] vdd 0.63fF
C983 la_data_out[18] vdd 0.63fF
C984 la_data_in[18] vdd 0.63fF
C985 la_oenb[17] vdd 0.63fF
C986 la_data_out[17] vdd 0.63fF
C987 la_data_in[17] vdd 0.63fF
C988 la_oenb[16] vdd 0.63fF
C989 la_data_out[16] vdd 0.63fF
C990 la_data_in[16] vdd 0.63fF
C991 la_oenb[15] vdd 0.63fF
C992 la_data_out[15] vdd 0.63fF
C993 la_data_in[15] vdd 0.63fF
C994 la_oenb[14] vdd 0.63fF
C995 la_data_out[14] vdd 0.63fF
C996 la_data_in[14] vdd 0.63fF
C997 la_oenb[13] vdd 0.63fF
C998 la_data_out[13] vdd 0.63fF
C999 la_data_in[13] vdd 0.63fF
C1000 la_oenb[12] vdd 0.63fF
C1001 la_data_out[12] vdd 0.63fF
C1002 la_data_in[12] vdd 0.63fF
C1003 la_oenb[11] vdd 0.63fF
C1004 la_data_out[11] vdd 0.63fF
C1005 la_data_in[11] vdd 0.63fF
C1006 la_oenb[10] vdd 0.63fF
C1007 la_data_out[10] vdd 0.63fF
C1008 la_data_in[10] vdd 0.63fF
C1009 la_oenb[9] vdd 0.63fF
C1010 la_data_out[9] vdd 0.63fF
C1011 la_data_in[9] vdd 0.63fF
C1012 la_oenb[8] vdd 0.63fF
C1013 la_data_out[8] vdd 0.63fF
C1014 la_data_in[8] vdd 0.63fF
C1015 la_oenb[7] vdd 0.63fF
C1016 la_data_out[7] vdd 0.63fF
C1017 la_data_in[7] vdd 0.63fF
C1018 la_oenb[6] vdd 0.63fF
C1019 la_data_out[6] vdd 0.63fF
C1020 la_data_in[6] vdd 0.63fF
C1021 la_oenb[5] vdd 0.63fF
C1022 la_data_out[5] vdd 0.63fF
C1023 la_data_in[5] vdd 0.63fF
C1024 la_oenb[4] vdd 0.63fF
C1025 la_data_out[4] vdd 0.63fF
C1026 la_data_in[4] vdd 0.63fF
C1027 la_oenb[3] vdd 0.63fF
C1028 la_data_out[3] vdd 0.63fF
C1029 la_data_in[3] vdd 0.63fF
C1030 la_oenb[2] vdd 0.63fF
C1031 la_data_out[2] vdd 0.63fF
C1032 la_data_in[2] vdd 0.63fF
C1033 la_oenb[1] vdd 0.63fF
C1034 la_data_out[1] vdd 0.63fF
C1035 la_data_in[1] vdd 0.63fF
C1036 la_oenb[0] vdd 0.63fF
C1037 la_data_out[0] vdd 0.63fF
C1038 la_data_in[0] vdd 0.63fF
C1039 wbs_dat_o[31] vdd 0.63fF
C1040 wbs_dat_i[31] vdd 0.63fF
C1041 wbs_adr_i[31] vdd 0.63fF
C1042 wbs_dat_o[30] vdd 0.63fF
C1043 wbs_dat_i[30] vdd 0.63fF
C1044 wbs_adr_i[30] vdd 0.63fF
C1045 wbs_dat_o[29] vdd 0.63fF
C1046 wbs_dat_i[29] vdd 0.63fF
C1047 wbs_adr_i[29] vdd 0.63fF
C1048 wbs_dat_o[28] vdd 0.63fF
C1049 wbs_dat_i[28] vdd 0.63fF
C1050 wbs_adr_i[28] vdd 0.63fF
C1051 wbs_dat_o[27] vdd 0.63fF
C1052 wbs_dat_i[27] vdd 0.63fF
C1053 wbs_adr_i[27] vdd 0.63fF
C1054 wbs_dat_o[26] vdd 0.63fF
C1055 wbs_dat_i[26] vdd 0.63fF
C1056 wbs_adr_i[26] vdd 0.63fF
C1057 wbs_dat_o[25] vdd 0.63fF
C1058 wbs_dat_i[25] vdd 0.63fF
C1059 wbs_adr_i[25] vdd 0.63fF
C1060 wbs_dat_o[24] vdd 0.63fF
C1061 wbs_dat_i[24] vdd 0.63fF
C1062 wbs_adr_i[24] vdd 0.63fF
C1063 wbs_dat_o[23] vdd 0.63fF
C1064 wbs_dat_i[23] vdd 0.63fF
C1065 wbs_adr_i[23] vdd 0.63fF
C1066 wbs_dat_o[22] vdd 0.63fF
C1067 wbs_dat_i[22] vdd 0.63fF
C1068 wbs_adr_i[22] vdd 0.63fF
C1069 wbs_dat_o[21] vdd 0.63fF
C1070 wbs_dat_i[21] vdd 0.63fF
C1071 wbs_adr_i[21] vdd 0.63fF
C1072 wbs_dat_o[20] vdd 0.63fF
C1073 wbs_dat_i[20] vdd 0.63fF
C1074 wbs_adr_i[20] vdd 0.63fF
C1075 wbs_dat_o[19] vdd 0.63fF
C1076 wbs_dat_i[19] vdd 0.63fF
C1077 wbs_adr_i[19] vdd 0.63fF
C1078 wbs_dat_o[18] vdd 0.63fF
C1079 wbs_dat_i[18] vdd 0.63fF
C1080 wbs_adr_i[18] vdd 0.63fF
C1081 wbs_dat_o[17] vdd 0.63fF
C1082 wbs_dat_i[17] vdd 0.63fF
C1083 wbs_adr_i[17] vdd 0.63fF
C1084 wbs_dat_o[16] vdd 0.63fF
C1085 wbs_dat_i[16] vdd 0.63fF
C1086 wbs_adr_i[16] vdd 0.63fF
C1087 wbs_dat_o[15] vdd 0.63fF
C1088 wbs_dat_i[15] vdd 0.63fF
C1089 wbs_adr_i[15] vdd 0.63fF
C1090 wbs_dat_o[14] vdd 0.63fF
C1091 wbs_dat_i[14] vdd 0.63fF
C1092 wbs_adr_i[14] vdd 0.63fF
C1093 wbs_dat_o[13] vdd 0.63fF
C1094 wbs_dat_i[13] vdd 0.63fF
C1095 wbs_adr_i[13] vdd 0.63fF
C1096 wbs_dat_o[12] vdd 0.63fF
C1097 wbs_dat_i[12] vdd 0.63fF
C1098 wbs_adr_i[12] vdd 0.63fF
C1099 wbs_dat_o[11] vdd 0.63fF
C1100 wbs_dat_i[11] vdd 0.63fF
C1101 wbs_adr_i[11] vdd 0.63fF
C1102 wbs_dat_o[10] vdd 0.63fF
C1103 wbs_dat_i[10] vdd 0.63fF
C1104 wbs_adr_i[10] vdd 0.63fF
C1105 wbs_dat_o[9] vdd 0.63fF
C1106 wbs_dat_i[9] vdd 0.63fF
C1107 wbs_adr_i[9] vdd 0.63fF
C1108 wbs_dat_o[8] vdd 0.63fF
C1109 wbs_dat_i[8] vdd 0.63fF
C1110 wbs_adr_i[8] vdd 0.63fF
C1111 wbs_dat_o[7] vdd 0.63fF
C1112 wbs_dat_i[7] vdd 0.63fF
C1113 wbs_adr_i[7] vdd 0.63fF
C1114 wbs_dat_o[6] vdd 0.63fF
C1115 wbs_dat_i[6] vdd 0.63fF
C1116 wbs_adr_i[6] vdd 0.63fF
C1117 wbs_dat_o[5] vdd 0.63fF
C1118 wbs_dat_i[5] vdd 0.63fF
C1119 wbs_adr_i[5] vdd 0.63fF
C1120 wbs_dat_o[4] vdd 0.63fF
C1121 wbs_dat_i[4] vdd 0.63fF
C1122 wbs_adr_i[4] vdd 0.63fF
C1123 wbs_sel_i[3] vdd 0.63fF
C1124 wbs_dat_o[3] vdd 0.63fF
C1125 wbs_dat_i[3] vdd 0.63fF
C1126 wbs_adr_i[3] vdd 0.63fF
C1127 wbs_sel_i[2] vdd 0.63fF
C1128 wbs_dat_o[2] vdd 0.63fF
C1129 wbs_dat_i[2] vdd 0.63fF
C1130 wbs_adr_i[2] vdd 0.63fF
C1131 wbs_sel_i[1] vdd 0.63fF
C1132 wbs_dat_o[1] vdd 0.63fF
C1133 wbs_dat_i[1] vdd 0.63fF
C1134 wbs_adr_i[1] vdd 0.63fF
C1135 wbs_sel_i[0] vdd 0.63fF
C1136 wbs_dat_o[0] vdd 0.63fF
C1137 wbs_dat_i[0] vdd 0.63fF
C1138 wbs_adr_i[0] vdd 0.63fF
C1139 wbs_we_i vdd 0.63fF
C1140 wbs_stb_i vdd 0.63fF
C1141 wbs_cyc_i vdd 0.63fF
C1142 wbs_ack_o vdd 0.63fF
C1143 wb_rst_i vdd 0.63fF
C1144 wb_clk_i vdd 0.63fF
C1145 divider_0/and_0/Z1 vdd 0.32fF
C1146 divider_0/and_0/B vdd 2.06fF
C1147 divider_0/and_0/out1 vdd 1.27fF
C1148 divider_0/tspc_2/a_630_n680# vdd 0.53fF
C1149 divider_0/tspc_2/Z4 vdd 0.41fF
C1150 divider_0/Out vdd 0.70fF
C1151 divider_0/tspc_2/Z3 vdd 1.33fF
C1152 divider_0/tspc_2/Z2 vdd 0.91fF
C1153 divider_0/tspc_2/Z1 vdd 0.42fF
C1154 divider_0/tspc_1/Q vdd 1.46fF
C1155 divider_0/nor_1/B vdd 5.20fF
C1156 divider_0/tspc_1/a_630_n680# vdd 0.53fF
C1157 divider_0/tspc_1/Z4 vdd 0.41fF
C1158 divider_0/tspc_1/Z3 vdd 1.33fF
C1159 divider_0/tspc_1/Z2 vdd 0.91fF
C1160 divider_0/tspc_1/Z1 vdd 0.42fF
C1161 divider_0/tspc_0/Q vdd 1.95fF
C1162 divider_0/nor_0/B vdd 4.86fF
C1163 divider_0/tspc_0/a_630_n680# vdd 0.53fF
C1164 divider_0/tspc_0/Z4 vdd 0.41fF
C1165 divider_0/tspc_0/Z3 vdd 1.33fF
C1166 divider_0/tspc_0/Z2 vdd 0.91fF
C1167 divider_0/tspc_0/Z1 vdd 0.42fF
C1168 divider_0/nor_0/A vdd 4.47fF
C1169 divider_0/clk vdd 5.27fF
C1170 divider_0/prescaler_0/nand_1/z1 vdd 0.20fF
C1171 divider_0/prescaler_0/tspc_2/D vdd 2.15fF
C1172 divider_0/and_0/OUT vdd 3.38fF
C1173 divider_0/prescaler_0/nand_0/z1 vdd 0.20fF
C1174 divider_0/vdd vdd 23.71fF
C1175 divider_0/prescaler_0/tspc_1/Q vdd 1.91fF
C1176 divider_0/prescaler_0/tspc_2/Q vdd 2.54fF
C1177 divider_0/prescaler_0/tspc_2/a_630_n680# vdd 0.53fF
C1178 divider_0/prescaler_0/tspc_2/Z4 vdd 0.41fF
C1179 divider_0/prescaler_0/tspc_2/Z3 vdd 1.33fF
C1180 divider_0/prescaler_0/tspc_2/Z2 vdd 0.91fF
C1181 divider_0/prescaler_0/tspc_2/Z1 vdd 0.43fF
C1182 divider_0/prescaler_0/tspc_2/a_740_n680# vdd 1.37fF
C1183 divider_0/prescaler_0/tspc_1/a_630_n680# vdd 0.53fF
C1184 divider_0/prescaler_0/tspc_1/Z4 vdd 0.41fF
C1185 divider_0/prescaler_0/tspc_1/Z3 vdd 1.33fF
C1186 divider_0/prescaler_0/tspc_1/Z2 vdd 0.91fF
C1187 divider_0/prescaler_0/tspc_1/Z1 vdd 0.42fF
C1188 divider_0/prescaler_0/m1_2700_2190# vdd 3.36fF
C1189 divider_0/prescaler_0/tspc_0/a_630_n680# vdd 0.53fF
C1190 divider_0/gnd vdd 21.09fF
C1191 divider_0/prescaler_0/tspc_0/Z4 vdd 0.42fF
C1192 divider_0/prescaler_0/Out vdd 3.22fF
C1193 divider_0/prescaler_0/tspc_0/Z3 vdd 1.33fF
C1194 divider_0/prescaler_0/tspc_0/Z2 vdd 0.91fF
C1195 divider_0/prescaler_0/tspc_0/Z1 vdd 0.44fF
C1196 divider_0/prescaler_0/tspc_0/D vdd 1.79fF
C1197 divider_0/prescaler_0/tspc_0/a_740_n680# vdd 1.37fF
C1198 divider_0/nor_1/Z1 vdd 0.60fF
C1199 divider_0/mc2 vdd 3.52fF
C1200 divider_0/and_0/A vdd 1.65fF
C1201 divider_0/nor_0/Z1 vdd 0.60fF
C1202 ro_complete_0/cbank_2/switch_0/vin vdd 1.30fF
C1203 ro_complete_0/cbank_2/v vdd 15.52fF
C1204 ro_complete_0/cbank_2/switch_5/vin vdd 1.06fF
C1205 ro_complete_0/a5 vdd 5.32fF
C1206 ro_complete_0/cbank_2/switch_4/vin vdd 1.16fF
C1207 ro_complete_0/a4 vdd 5.44fF
C1208 ro_complete_0/cbank_2/switch_2/vin vdd 0.95fF
C1209 ro_complete_0/a2 vdd 5.61fF
C1210 ro_complete_0/cbank_2/switch_3/vin vdd 1.30fF
C1211 ro_complete_0/a3 vdd 7.09fF
C1212 ro_complete_0/cbank_2/switch_1/vin vdd 1.53fF
C1213 ro_complete_0/a1 vdd 5.46fF
C1214 ro_complete_0/a0 vdd 7.97fF
C1215 ro_complete_0/cbank_1/switch_0/vin vdd 1.30fF
C1216 ro_complete_0/cbank_1/v vdd 16.22fF
C1217 ro_complete_0/cbank_1/switch_5/vin vdd 1.06fF
C1218 ro_complete_0/cbank_1/switch_4/vin vdd 1.16fF
C1219 ro_complete_0/cbank_1/switch_2/vin vdd 0.95fF
C1220 ro_complete_0/cbank_1/switch_3/vin vdd 1.30fF
C1221 ro_complete_0/cbank_1/switch_1/vin vdd 1.53fF
C1222 ro_complete_0/cbank_0/switch_0/vin vdd 1.30fF
C1223 ro_complete_0/cbank_0/v vdd 14.76fF
C1224 ro_complete_0/cbank_0/switch_5/vin vdd 1.06fF
C1225 ro_complete_0/cbank_0/switch_4/vin vdd 1.16fF
C1226 ro_complete_0/cbank_0/switch_2/vin vdd 0.95fF
C1227 ro_complete_0/cbank_0/switch_3/vin vdd 1.30fF
C1228 ro_complete_0/cbank_0/switch_1/vin vdd 1.53fF
C1229 ro_complete_0/ro_var_extend_0/vcont vdd 0.46fF **FLOATING
C1230 cp_0/a_7110_n2840# vdd 0.17fF
C1231 cp_0/a_3060_n2840# vdd 1.71fF
C1232 cp_0/down vdd 0.90fF
C1233 cp_0/vbias vdd 2.41fF
C1234 cp_0/a_7110_0# vdd 0.17fF
C1235 cp_0/a_3060_0# vdd 1.65fF
C1236 cp_0/a_1710_0# vdd 5.76fF
C1237 cp_0/upbar vdd 0.88fF
C1238 cp_0/out vdd 5.14fF
C1239 cp_0/a_1710_n2840# vdd 4.85fF
C1240 cp_0/a_10_n50# vdd 2.96fF
C1241 pd_0/and_pd_0/Z1 vdd 0.20fF
C1242 pd_0/and_pd_0/Out1 vdd 2.01fF
C1243 pd_0/tspc_r_1/z5 vdd 0.53fF
C1244 pd_0/tspc_r_1/Z4 vdd 0.53fF
C1245 pd_0/R vdd 2.48fF
C1246 pd_0/tspc_r_1/Qbar vdd 0.61fF
C1247 pd_0/tspc_r_1/Z2 vdd 1.05fF
C1248 pd_0/tspc_r_1/Z1 vdd 0.66fF
C1249 pd_0/DOWN vdd 2.21fF
C1250 pd_0/tspc_r_1/Qbar1 vdd 1.17fF
C1251 pd_0/tspc_r_1/Z3 vdd 1.79fF
C1252 pd_0/DIV vdd 1.78fF
C1253 pd_0/tspc_r_0/z5 vdd 0.53fF
C1254 pd_0/tspc_r_0/Z4 vdd 0.53fF
C1255 GND vdd 7.48fF
C1256 pd_0/tspc_r_0/Qbar vdd 0.69fF
C1257 pd_0/tspc_r_0/Z2 vdd 1.07fF
C1258 pd_0/tspc_r_0/Z1 vdd 0.66fF
C1259 pd_0/UP vdd 2.15fF
C1260 pd_0/tspc_r_0/Qbar1 vdd 1.17fF
C1261 pd_0/tspc_r_0/Z3 vdd 1.79fF
C1262 pd_0/REF vdd 1.76fF
.ends
