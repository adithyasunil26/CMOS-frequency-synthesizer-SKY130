magic
tech sky130A
timestamp 1640906950
<< nwell >>
rect -245 1860 4500 2030
rect -245 -80 4495 1860
<< nmos >>
rect 5 -1420 185 -520
rect 675 -1420 855 -520
rect 1350 -1420 1530 -520
rect 2025 -1420 2205 -520
rect 2700 -1420 2880 -520
rect 3375 -1420 3555 -520
rect 4050 -1420 4230 -520
<< pmos >>
rect 5 0 185 1800
rect 675 0 855 1800
rect 1350 0 1530 1800
rect 2025 0 2205 1800
rect 2700 0 2880 1800
rect 3375 0 3555 1800
rect 4050 0 4230 1800
<< ndiff >>
rect -185 -600 5 -520
rect -185 -700 -140 -600
rect -40 -700 5 -600
rect -185 -810 5 -700
rect -185 -910 -140 -810
rect -40 -910 5 -810
rect -185 -1020 5 -910
rect -185 -1120 -140 -1020
rect -40 -1120 5 -1020
rect -185 -1230 5 -1120
rect -185 -1330 -140 -1230
rect -40 -1330 5 -1230
rect -185 -1420 5 -1330
rect 185 -600 375 -520
rect 185 -700 230 -600
rect 330 -700 375 -600
rect 185 -810 375 -700
rect 185 -910 230 -810
rect 330 -910 375 -810
rect 185 -1020 375 -910
rect 185 -1120 230 -1020
rect 330 -1120 375 -1020
rect 185 -1230 375 -1120
rect 185 -1330 230 -1230
rect 330 -1330 375 -1230
rect 185 -1420 375 -1330
rect 485 -600 675 -520
rect 485 -700 530 -600
rect 630 -700 675 -600
rect 485 -810 675 -700
rect 485 -910 530 -810
rect 630 -910 675 -810
rect 485 -1020 675 -910
rect 485 -1120 530 -1020
rect 630 -1120 675 -1020
rect 485 -1230 675 -1120
rect 485 -1330 530 -1230
rect 630 -1330 675 -1230
rect 485 -1415 675 -1330
rect 515 -1420 675 -1415
rect 855 -600 1045 -520
rect 855 -700 900 -600
rect 1000 -700 1045 -600
rect 855 -810 1045 -700
rect 855 -910 900 -810
rect 1000 -910 1045 -810
rect 855 -1020 1045 -910
rect 855 -1120 900 -1020
rect 1000 -1120 1045 -1020
rect 855 -1230 1045 -1120
rect 855 -1330 900 -1230
rect 1000 -1330 1045 -1230
rect 855 -1420 1045 -1330
rect 1160 -600 1350 -520
rect 1160 -700 1205 -600
rect 1305 -700 1350 -600
rect 1160 -810 1350 -700
rect 1160 -910 1205 -810
rect 1305 -910 1350 -810
rect 1160 -1020 1350 -910
rect 1160 -1120 1205 -1020
rect 1305 -1120 1350 -1020
rect 1160 -1230 1350 -1120
rect 1160 -1330 1205 -1230
rect 1305 -1330 1350 -1230
rect 1160 -1420 1350 -1330
rect 1530 -600 1720 -520
rect 1530 -700 1575 -600
rect 1675 -700 1720 -600
rect 1530 -810 1720 -700
rect 1530 -910 1575 -810
rect 1675 -910 1720 -810
rect 1530 -1020 1720 -910
rect 1530 -1120 1575 -1020
rect 1675 -1120 1720 -1020
rect 1530 -1230 1720 -1120
rect 1530 -1330 1575 -1230
rect 1675 -1330 1720 -1230
rect 1530 -1420 1720 -1330
rect 1835 -600 2025 -520
rect 1835 -700 1880 -600
rect 1980 -700 2025 -600
rect 1835 -810 2025 -700
rect 1835 -910 1880 -810
rect 1980 -910 2025 -810
rect 1835 -1020 2025 -910
rect 1835 -1120 1880 -1020
rect 1980 -1120 2025 -1020
rect 1835 -1230 2025 -1120
rect 1835 -1330 1880 -1230
rect 1980 -1330 2025 -1230
rect 1835 -1420 2025 -1330
rect 2205 -600 2395 -520
rect 2205 -700 2250 -600
rect 2350 -700 2395 -600
rect 2205 -810 2395 -700
rect 2205 -910 2250 -810
rect 2350 -910 2395 -810
rect 2205 -1020 2395 -910
rect 2205 -1120 2250 -1020
rect 2350 -1120 2395 -1020
rect 2205 -1230 2395 -1120
rect 2205 -1330 2250 -1230
rect 2350 -1330 2395 -1230
rect 2205 -1420 2395 -1330
rect 2510 -600 2700 -520
rect 2510 -700 2555 -600
rect 2655 -700 2700 -600
rect 2510 -810 2700 -700
rect 2510 -910 2555 -810
rect 2655 -910 2700 -810
rect 2510 -1020 2700 -910
rect 2510 -1120 2555 -1020
rect 2655 -1120 2700 -1020
rect 2510 -1230 2700 -1120
rect 2510 -1330 2555 -1230
rect 2655 -1330 2700 -1230
rect 2510 -1420 2700 -1330
rect 2880 -600 3070 -520
rect 2880 -700 2925 -600
rect 3025 -700 3070 -600
rect 2880 -810 3070 -700
rect 2880 -910 2925 -810
rect 3025 -910 3070 -810
rect 2880 -1020 3070 -910
rect 2880 -1120 2925 -1020
rect 3025 -1120 3070 -1020
rect 2880 -1230 3070 -1120
rect 2880 -1330 2925 -1230
rect 3025 -1330 3070 -1230
rect 2880 -1420 3070 -1330
rect 3185 -600 3375 -520
rect 3185 -700 3230 -600
rect 3330 -700 3375 -600
rect 3185 -810 3375 -700
rect 3185 -910 3230 -810
rect 3330 -910 3375 -810
rect 3185 -1020 3375 -910
rect 3185 -1120 3230 -1020
rect 3330 -1120 3375 -1020
rect 3185 -1230 3375 -1120
rect 3185 -1330 3230 -1230
rect 3330 -1330 3375 -1230
rect 3185 -1420 3375 -1330
rect 3555 -600 3745 -520
rect 3555 -700 3600 -600
rect 3700 -700 3745 -600
rect 3555 -810 3745 -700
rect 3555 -910 3600 -810
rect 3700 -910 3745 -810
rect 3555 -1020 3745 -910
rect 3555 -1120 3600 -1020
rect 3700 -1120 3745 -1020
rect 3555 -1230 3745 -1120
rect 3555 -1330 3600 -1230
rect 3700 -1330 3745 -1230
rect 3555 -1420 3745 -1330
rect 3860 -600 4050 -520
rect 3860 -700 3905 -600
rect 4005 -700 4050 -600
rect 3860 -810 4050 -700
rect 3860 -910 3905 -810
rect 4005 -910 4050 -810
rect 3860 -1020 4050 -910
rect 3860 -1120 3905 -1020
rect 4005 -1120 4050 -1020
rect 3860 -1230 4050 -1120
rect 3860 -1330 3905 -1230
rect 4005 -1330 4050 -1230
rect 3860 -1420 4050 -1330
rect 4230 -600 4420 -520
rect 4230 -700 4275 -600
rect 4375 -700 4420 -600
rect 4230 -810 4420 -700
rect 4230 -910 4275 -810
rect 4375 -910 4420 -810
rect 4230 -1020 4420 -910
rect 4230 -1120 4275 -1020
rect 4375 -1120 4420 -1020
rect 4230 -1230 4420 -1120
rect 4230 -1330 4275 -1230
rect 4375 -1330 4420 -1230
rect 4230 -1420 4420 -1330
<< pdiff >>
rect -185 1715 5 1800
rect -185 1615 -140 1715
rect -40 1615 5 1715
rect -185 1430 5 1615
rect -185 1330 -140 1430
rect -40 1330 5 1430
rect -185 1115 5 1330
rect -185 1015 -140 1115
rect -40 1015 5 1115
rect -185 800 5 1015
rect -185 700 -140 800
rect -40 700 5 800
rect -185 465 5 700
rect -185 365 -140 465
rect -40 365 5 465
rect -185 140 5 365
rect -185 40 -140 140
rect -40 40 5 140
rect -185 0 5 40
rect 185 1715 375 1800
rect 185 1615 230 1715
rect 330 1615 375 1715
rect 185 1430 375 1615
rect 185 1330 230 1430
rect 330 1330 375 1430
rect 185 1115 375 1330
rect 185 1015 230 1115
rect 330 1015 375 1115
rect 185 800 375 1015
rect 185 700 230 800
rect 330 700 375 800
rect 185 465 375 700
rect 185 365 230 465
rect 330 365 375 465
rect 185 140 375 365
rect 185 40 230 140
rect 330 40 375 140
rect 185 0 375 40
rect 485 1715 675 1800
rect 485 1615 530 1715
rect 630 1615 675 1715
rect 485 1430 675 1615
rect 485 1330 530 1430
rect 630 1330 675 1430
rect 485 1115 675 1330
rect 485 1015 530 1115
rect 630 1015 675 1115
rect 485 800 675 1015
rect 485 700 530 800
rect 630 700 675 800
rect 485 465 675 700
rect 485 365 530 465
rect 630 365 675 465
rect 485 140 675 365
rect 485 40 530 140
rect 630 40 675 140
rect 485 0 675 40
rect 855 1715 1045 1800
rect 855 1615 900 1715
rect 1000 1615 1045 1715
rect 855 1430 1045 1615
rect 855 1330 900 1430
rect 1000 1330 1045 1430
rect 855 1115 1045 1330
rect 855 1015 900 1115
rect 1000 1015 1045 1115
rect 855 800 1045 1015
rect 855 700 900 800
rect 1000 700 1045 800
rect 855 465 1045 700
rect 855 365 900 465
rect 1000 365 1045 465
rect 855 140 1045 365
rect 855 40 900 140
rect 1000 40 1045 140
rect 855 0 1045 40
rect 1160 1715 1350 1800
rect 1160 1615 1205 1715
rect 1305 1615 1350 1715
rect 1160 1430 1350 1615
rect 1160 1330 1205 1430
rect 1305 1330 1350 1430
rect 1160 1115 1350 1330
rect 1160 1015 1205 1115
rect 1305 1015 1350 1115
rect 1160 800 1350 1015
rect 1160 700 1205 800
rect 1305 700 1350 800
rect 1160 465 1350 700
rect 1160 365 1205 465
rect 1305 365 1350 465
rect 1160 140 1350 365
rect 1160 40 1205 140
rect 1305 40 1350 140
rect 1160 0 1350 40
rect 1530 1715 1720 1800
rect 1530 1615 1575 1715
rect 1675 1615 1720 1715
rect 1530 1430 1720 1615
rect 1530 1330 1575 1430
rect 1675 1330 1720 1430
rect 1530 1115 1720 1330
rect 1530 1015 1575 1115
rect 1675 1015 1720 1115
rect 1530 800 1720 1015
rect 1530 700 1575 800
rect 1675 700 1720 800
rect 1530 465 1720 700
rect 1530 365 1575 465
rect 1675 365 1720 465
rect 1530 145 1720 365
rect 1530 45 1575 145
rect 1675 45 1720 145
rect 1530 0 1720 45
rect 1835 1715 2025 1800
rect 1835 1615 1880 1715
rect 1980 1615 2025 1715
rect 1835 1430 2025 1615
rect 1835 1330 1880 1430
rect 1980 1330 2025 1430
rect 1835 1115 2025 1330
rect 1835 1015 1880 1115
rect 1980 1015 2025 1115
rect 1835 800 2025 1015
rect 1835 700 1880 800
rect 1980 700 2025 800
rect 1835 465 2025 700
rect 1835 365 1880 465
rect 1980 365 2025 465
rect 1835 145 2025 365
rect 1835 45 1880 145
rect 1980 45 2025 145
rect 1835 0 2025 45
rect 2205 1715 2395 1800
rect 2205 1615 2250 1715
rect 2350 1615 2395 1715
rect 2205 1430 2395 1615
rect 2205 1330 2250 1430
rect 2350 1330 2395 1430
rect 2205 1115 2395 1330
rect 2205 1015 2250 1115
rect 2350 1015 2395 1115
rect 2205 800 2395 1015
rect 2205 700 2250 800
rect 2350 700 2395 800
rect 2205 465 2395 700
rect 2205 365 2250 465
rect 2350 365 2395 465
rect 2205 145 2395 365
rect 2205 45 2250 145
rect 2350 45 2395 145
rect 2205 0 2395 45
rect 2510 1715 2700 1800
rect 2510 1615 2555 1715
rect 2655 1615 2700 1715
rect 2510 1430 2700 1615
rect 2510 1330 2555 1430
rect 2655 1330 2700 1430
rect 2510 1115 2700 1330
rect 2510 1015 2555 1115
rect 2655 1015 2700 1115
rect 2510 800 2700 1015
rect 2510 700 2555 800
rect 2655 700 2700 800
rect 2510 465 2700 700
rect 2510 365 2555 465
rect 2655 365 2700 465
rect 2510 145 2700 365
rect 2510 45 2555 145
rect 2655 45 2700 145
rect 2510 0 2700 45
rect 2880 1715 3070 1800
rect 2880 1615 2925 1715
rect 3025 1615 3070 1715
rect 2880 1430 3070 1615
rect 2880 1330 2925 1430
rect 3025 1330 3070 1430
rect 2880 1115 3070 1330
rect 2880 1015 2925 1115
rect 3025 1015 3070 1115
rect 2880 800 3070 1015
rect 2880 700 2925 800
rect 3025 700 3070 800
rect 2880 465 3070 700
rect 2880 365 2925 465
rect 3025 365 3070 465
rect 2880 140 3070 365
rect 2880 40 2925 140
rect 3025 40 3070 140
rect 2880 0 3070 40
rect 3185 1715 3375 1800
rect 3185 1615 3230 1715
rect 3330 1615 3375 1715
rect 3185 1430 3375 1615
rect 3185 1330 3230 1430
rect 3330 1330 3375 1430
rect 3185 1115 3375 1330
rect 3185 1015 3230 1115
rect 3330 1015 3375 1115
rect 3185 800 3375 1015
rect 3185 700 3230 800
rect 3330 700 3375 800
rect 3185 465 3375 700
rect 3185 365 3230 465
rect 3330 365 3375 465
rect 3185 140 3375 365
rect 3185 40 3230 140
rect 3330 40 3375 140
rect 3185 0 3375 40
rect 3555 1715 3745 1800
rect 3555 1615 3600 1715
rect 3700 1615 3745 1715
rect 3555 1430 3745 1615
rect 3555 1330 3600 1430
rect 3700 1330 3745 1430
rect 3555 1115 3745 1330
rect 3555 1015 3600 1115
rect 3700 1015 3745 1115
rect 3555 800 3745 1015
rect 3555 700 3600 800
rect 3700 700 3745 800
rect 3555 465 3745 700
rect 3555 365 3600 465
rect 3700 365 3745 465
rect 3555 140 3745 365
rect 3555 40 3600 140
rect 3700 40 3745 140
rect 3555 0 3745 40
rect 3860 1715 4050 1800
rect 3860 1615 3905 1715
rect 4005 1615 4050 1715
rect 3860 1430 4050 1615
rect 3860 1330 3905 1430
rect 4005 1330 4050 1430
rect 3860 1115 4050 1330
rect 3860 1015 3905 1115
rect 4005 1015 4050 1115
rect 3860 800 4050 1015
rect 3860 700 3905 800
rect 4005 700 4050 800
rect 3860 465 4050 700
rect 3860 365 3905 465
rect 4005 365 4050 465
rect 3860 140 4050 365
rect 3860 40 3905 140
rect 4005 40 4050 140
rect 3860 0 4050 40
rect 4230 1715 4420 1800
rect 4230 1615 4275 1715
rect 4375 1615 4420 1715
rect 4230 1430 4420 1615
rect 4230 1330 4275 1430
rect 4375 1330 4420 1430
rect 4230 1115 4420 1330
rect 4230 1015 4275 1115
rect 4375 1015 4420 1115
rect 4230 800 4420 1015
rect 4230 700 4275 800
rect 4375 700 4420 800
rect 4230 465 4420 700
rect 4230 365 4275 465
rect 4375 365 4420 465
rect 4230 140 4420 365
rect 4230 40 4275 140
rect 4375 40 4420 140
rect 4230 0 4420 40
<< ndiffc >>
rect -140 -700 -40 -600
rect -140 -910 -40 -810
rect -140 -1120 -40 -1020
rect -140 -1330 -40 -1230
rect 230 -700 330 -600
rect 230 -910 330 -810
rect 230 -1120 330 -1020
rect 230 -1330 330 -1230
rect 530 -700 630 -600
rect 530 -910 630 -810
rect 530 -1120 630 -1020
rect 530 -1330 630 -1230
rect 900 -700 1000 -600
rect 900 -910 1000 -810
rect 900 -1120 1000 -1020
rect 900 -1330 1000 -1230
rect 1205 -700 1305 -600
rect 1205 -910 1305 -810
rect 1205 -1120 1305 -1020
rect 1205 -1330 1305 -1230
rect 1575 -700 1675 -600
rect 1575 -910 1675 -810
rect 1575 -1120 1675 -1020
rect 1575 -1330 1675 -1230
rect 1880 -700 1980 -600
rect 1880 -910 1980 -810
rect 1880 -1120 1980 -1020
rect 1880 -1330 1980 -1230
rect 2250 -700 2350 -600
rect 2250 -910 2350 -810
rect 2250 -1120 2350 -1020
rect 2250 -1330 2350 -1230
rect 2555 -700 2655 -600
rect 2555 -910 2655 -810
rect 2555 -1120 2655 -1020
rect 2555 -1330 2655 -1230
rect 2925 -700 3025 -600
rect 2925 -910 3025 -810
rect 2925 -1120 3025 -1020
rect 2925 -1330 3025 -1230
rect 3230 -700 3330 -600
rect 3230 -910 3330 -810
rect 3230 -1120 3330 -1020
rect 3230 -1330 3330 -1230
rect 3600 -700 3700 -600
rect 3600 -910 3700 -810
rect 3600 -1120 3700 -1020
rect 3600 -1330 3700 -1230
rect 3905 -700 4005 -600
rect 3905 -910 4005 -810
rect 3905 -1120 4005 -1020
rect 3905 -1330 4005 -1230
rect 4275 -700 4375 -600
rect 4275 -910 4375 -810
rect 4275 -1120 4375 -1020
rect 4275 -1330 4375 -1230
<< pdiffc >>
rect -140 1615 -40 1715
rect -140 1330 -40 1430
rect -140 1015 -40 1115
rect -140 700 -40 800
rect -140 365 -40 465
rect -140 40 -40 140
rect 230 1615 330 1715
rect 230 1330 330 1430
rect 230 1015 330 1115
rect 230 700 330 800
rect 230 365 330 465
rect 230 40 330 140
rect 530 1615 630 1715
rect 530 1330 630 1430
rect 530 1015 630 1115
rect 530 700 630 800
rect 530 365 630 465
rect 530 40 630 140
rect 900 1615 1000 1715
rect 900 1330 1000 1430
rect 900 1015 1000 1115
rect 900 700 1000 800
rect 900 365 1000 465
rect 900 40 1000 140
rect 1205 1615 1305 1715
rect 1205 1330 1305 1430
rect 1205 1015 1305 1115
rect 1205 700 1305 800
rect 1205 365 1305 465
rect 1205 40 1305 140
rect 1575 1615 1675 1715
rect 1575 1330 1675 1430
rect 1575 1015 1675 1115
rect 1575 700 1675 800
rect 1575 365 1675 465
rect 1575 45 1675 145
rect 1880 1615 1980 1715
rect 1880 1330 1980 1430
rect 1880 1015 1980 1115
rect 1880 700 1980 800
rect 1880 365 1980 465
rect 1880 45 1980 145
rect 2250 1615 2350 1715
rect 2250 1330 2350 1430
rect 2250 1015 2350 1115
rect 2250 700 2350 800
rect 2250 365 2350 465
rect 2250 45 2350 145
rect 2555 1615 2655 1715
rect 2555 1330 2655 1430
rect 2555 1015 2655 1115
rect 2555 700 2655 800
rect 2555 365 2655 465
rect 2555 45 2655 145
rect 2925 1615 3025 1715
rect 2925 1330 3025 1430
rect 2925 1015 3025 1115
rect 2925 700 3025 800
rect 2925 365 3025 465
rect 2925 40 3025 140
rect 3230 1615 3330 1715
rect 3230 1330 3330 1430
rect 3230 1015 3330 1115
rect 3230 700 3330 800
rect 3230 365 3330 465
rect 3230 40 3330 140
rect 3600 1615 3700 1715
rect 3600 1330 3700 1430
rect 3600 1015 3700 1115
rect 3600 700 3700 800
rect 3600 365 3700 465
rect 3600 40 3700 140
rect 3905 1615 4005 1715
rect 3905 1330 4005 1430
rect 3905 1015 4005 1115
rect 3905 700 4005 800
rect 3905 365 4005 465
rect 3905 40 4005 140
rect 4275 1615 4375 1715
rect 4275 1330 4375 1430
rect 4275 1015 4375 1115
rect 4275 700 4375 800
rect 4275 365 4375 465
rect 4275 40 4375 140
<< psubdiff >>
rect 2045 -1540 2190 -1525
rect 2045 -1650 2060 -1540
rect 2175 -1650 2190 -1540
rect 2045 -1665 2190 -1650
<< nsubdiff >>
rect 2045 1995 2190 2010
rect 2045 1885 2060 1995
rect 2175 1885 2190 1995
rect 2045 1875 2190 1885
<< psubdiffcont >>
rect 2060 -1650 2175 -1540
<< nsubdiffcont >>
rect 2060 1885 2175 1995
<< poly >>
rect 3405 1935 3525 1940
rect 3405 1835 3415 1935
rect 3515 1835 3525 1935
rect 3405 1825 3525 1835
rect 5 1800 185 1825
rect 675 1800 855 1825
rect 1350 1800 1530 1825
rect 2025 1800 2205 1825
rect 2700 1800 2880 1825
rect 3375 1800 3555 1825
rect 4050 1800 4230 1825
rect 5 -25 185 0
rect 675 -25 855 0
rect 1350 -25 1530 0
rect 2025 -25 2205 0
rect 2700 -25 2880 0
rect 3375 -25 3555 0
rect 4050 -25 4230 0
rect 40 -35 160 -25
rect 40 -135 50 -35
rect 150 -135 160 -35
rect 40 -145 160 -135
rect 705 -35 825 -25
rect 705 -135 715 -35
rect 815 -135 825 -35
rect 705 -145 825 -135
rect 1380 -35 1500 -25
rect 1380 -135 1390 -35
rect 1490 -135 1500 -35
rect 1380 -145 1500 -135
rect 2055 -35 2175 -25
rect 2055 -135 2065 -35
rect 2165 -135 2175 -35
rect 2055 -145 2175 -135
rect 2730 -35 2850 -25
rect 2730 -135 2740 -35
rect 2840 -135 2850 -35
rect 2730 -145 2850 -135
rect 3405 -35 3525 -25
rect 3405 -135 3415 -35
rect 3515 -135 3525 -35
rect 3405 -145 3525 -135
rect 4080 -35 4200 -25
rect 4080 -135 4090 -35
rect 4190 -135 4200 -35
rect 4080 -145 4200 -135
rect 40 -385 160 -375
rect 40 -485 50 -385
rect 150 -485 160 -385
rect 40 -495 160 -485
rect 705 -385 825 -375
rect 705 -485 715 -385
rect 815 -485 825 -385
rect 705 -495 825 -485
rect 1380 -385 1500 -375
rect 1380 -485 1390 -385
rect 1490 -485 1500 -385
rect 1380 -495 1500 -485
rect 2055 -385 2175 -375
rect 2055 -485 2065 -385
rect 2165 -485 2175 -385
rect 2055 -495 2175 -485
rect 2730 -385 2850 -375
rect 2730 -485 2740 -385
rect 2840 -485 2850 -385
rect 2730 -495 2850 -485
rect 3405 -385 3525 -375
rect 3405 -485 3415 -385
rect 3515 -485 3525 -385
rect 3405 -495 3525 -485
rect 4080 -385 4200 -375
rect 4080 -485 4090 -385
rect 4190 -485 4200 -385
rect 4080 -495 4200 -485
rect 5 -520 185 -495
rect 675 -520 855 -495
rect 1350 -520 1530 -495
rect 2025 -520 2205 -495
rect 2700 -520 2880 -495
rect 3375 -520 3555 -495
rect 4050 -520 4230 -495
rect 5 -1450 185 -1420
rect 675 -1450 855 -1420
rect 1350 -1450 1530 -1420
rect 2025 -1450 2205 -1420
rect 2700 -1450 2880 -1420
rect 3375 -1450 3555 -1420
rect 4050 -1450 4230 -1420
rect 3405 -1460 3525 -1450
rect 3405 -1560 3415 -1460
rect 3515 -1560 3525 -1460
rect 3405 -1570 3525 -1560
<< polycont >>
rect 3415 1835 3515 1935
rect 50 -135 150 -35
rect 715 -135 815 -35
rect 1390 -135 1490 -35
rect 2065 -135 2165 -35
rect 2740 -135 2840 -35
rect 3415 -135 3515 -35
rect 4090 -135 4190 -35
rect 50 -485 150 -385
rect 715 -485 815 -385
rect 1390 -485 1490 -385
rect 2065 -485 2165 -385
rect 2740 -485 2840 -385
rect 3415 -485 3515 -385
rect 4090 -485 4190 -385
rect 3415 -1560 3515 -1460
<< locali >>
rect -155 2000 -20 2010
rect -155 1890 -145 2000
rect -30 1890 -20 2000
rect -155 1785 -20 1890
rect 515 2000 650 2010
rect 515 1890 525 2000
rect 640 1890 650 2000
rect 515 1785 650 1890
rect 2050 1995 2185 2005
rect 2050 1885 2060 1995
rect 2175 1885 2185 1995
rect 2050 1880 2185 1885
rect 2905 2000 3040 2010
rect 2905 1890 2915 2000
rect 3030 1890 3040 2000
rect 2905 1785 3040 1890
rect 3405 1935 3525 1940
rect 3405 1835 3415 1935
rect 3515 1835 3525 1935
rect 3405 1825 3525 1835
rect -170 1715 -10 1785
rect -170 1615 -140 1715
rect -40 1615 -10 1715
rect -170 1430 -10 1615
rect -170 1330 -140 1430
rect -40 1330 -10 1430
rect -170 1115 -10 1330
rect -170 1015 -140 1115
rect -40 1015 -10 1115
rect -170 800 -10 1015
rect -170 700 -140 800
rect -40 700 -10 800
rect -170 465 -10 700
rect -170 365 -140 465
rect -40 365 -10 465
rect -170 140 -10 365
rect -170 40 -140 140
rect -40 40 -10 140
rect -170 15 -10 40
rect 200 1715 360 1785
rect 200 1615 230 1715
rect 330 1615 360 1715
rect 200 1430 360 1615
rect 200 1330 230 1430
rect 330 1330 360 1430
rect 200 1115 360 1330
rect 200 1015 230 1115
rect 330 1015 360 1115
rect 200 800 360 1015
rect 200 700 230 800
rect 330 700 360 800
rect 200 465 360 700
rect 200 365 230 465
rect 330 365 360 465
rect 200 140 360 365
rect 200 40 230 140
rect 330 40 360 140
rect 200 15 360 40
rect 500 1715 660 1785
rect 500 1615 530 1715
rect 630 1615 660 1715
rect 500 1430 660 1615
rect 500 1330 530 1430
rect 630 1330 660 1430
rect 500 1115 660 1330
rect 500 1015 530 1115
rect 630 1015 660 1115
rect 500 800 660 1015
rect 500 700 530 800
rect 630 700 660 800
rect 500 465 660 700
rect 500 365 530 465
rect 630 365 660 465
rect 500 140 660 365
rect 500 40 530 140
rect 630 40 660 140
rect 500 15 660 40
rect 870 1715 1030 1785
rect 870 1615 900 1715
rect 1000 1615 1030 1715
rect 870 1430 1030 1615
rect 870 1330 900 1430
rect 1000 1330 1030 1430
rect 870 1115 1030 1330
rect 870 1015 900 1115
rect 1000 1015 1030 1115
rect 870 800 1030 1015
rect 870 700 900 800
rect 1000 700 1030 800
rect 870 465 1030 700
rect 870 365 900 465
rect 1000 365 1030 465
rect 870 140 1030 365
rect 870 40 900 140
rect 1000 40 1030 140
rect 870 15 1030 40
rect 1175 1715 1335 1785
rect 1175 1615 1205 1715
rect 1305 1615 1335 1715
rect 1175 1430 1335 1615
rect 1175 1330 1205 1430
rect 1305 1330 1335 1430
rect 1175 1115 1335 1330
rect 1175 1015 1205 1115
rect 1305 1015 1335 1115
rect 1175 800 1335 1015
rect 1175 700 1205 800
rect 1305 700 1335 800
rect 1175 465 1335 700
rect 1175 365 1205 465
rect 1305 365 1335 465
rect 1175 140 1335 365
rect 1175 40 1205 140
rect 1305 40 1335 140
rect 1175 15 1335 40
rect 1545 1715 1705 1785
rect 1545 1615 1575 1715
rect 1675 1615 1705 1715
rect 1545 1430 1705 1615
rect 1545 1330 1575 1430
rect 1675 1330 1705 1430
rect 1545 1115 1705 1330
rect 1545 1015 1575 1115
rect 1675 1015 1705 1115
rect 1545 800 1705 1015
rect 1545 700 1575 800
rect 1675 700 1705 800
rect 1545 465 1705 700
rect 1545 365 1575 465
rect 1675 365 1705 465
rect 1545 145 1705 365
rect 1545 45 1575 145
rect 1675 45 1705 145
rect 1545 15 1705 45
rect 1850 1715 2010 1785
rect 1850 1615 1880 1715
rect 1980 1615 2010 1715
rect 1850 1430 2010 1615
rect 1850 1330 1880 1430
rect 1980 1330 2010 1430
rect 1850 1115 2010 1330
rect 1850 1015 1880 1115
rect 1980 1015 2010 1115
rect 1850 800 2010 1015
rect 1850 700 1880 800
rect 1980 700 2010 800
rect 1850 465 2010 700
rect 1850 365 1880 465
rect 1980 365 2010 465
rect 1850 145 2010 365
rect 1850 45 1880 145
rect 1980 45 2010 145
rect 1850 15 2010 45
rect 2220 1715 2380 1785
rect 2220 1615 2250 1715
rect 2350 1615 2380 1715
rect 2220 1430 2380 1615
rect 2220 1330 2250 1430
rect 2350 1330 2380 1430
rect 2220 1115 2380 1330
rect 2220 1015 2250 1115
rect 2350 1015 2380 1115
rect 2220 800 2380 1015
rect 2220 700 2250 800
rect 2350 700 2380 800
rect 2220 465 2380 700
rect 2220 365 2250 465
rect 2350 365 2380 465
rect 2220 145 2380 365
rect 2220 45 2250 145
rect 2350 45 2380 145
rect 2220 15 2380 45
rect 2525 1715 2685 1785
rect 2525 1615 2555 1715
rect 2655 1615 2685 1715
rect 2525 1430 2685 1615
rect 2525 1330 2555 1430
rect 2655 1330 2685 1430
rect 2525 1115 2685 1330
rect 2525 1015 2555 1115
rect 2655 1015 2685 1115
rect 2525 800 2685 1015
rect 2525 700 2555 800
rect 2655 700 2685 800
rect 2525 465 2685 700
rect 2525 365 2555 465
rect 2655 365 2685 465
rect 2525 145 2685 365
rect 2525 45 2555 145
rect 2655 45 2685 145
rect 2525 15 2685 45
rect 2895 1715 3055 1785
rect 2895 1615 2925 1715
rect 3025 1615 3055 1715
rect 2895 1430 3055 1615
rect 2895 1330 2925 1430
rect 3025 1330 3055 1430
rect 2895 1115 3055 1330
rect 2895 1015 2925 1115
rect 3025 1015 3055 1115
rect 2895 800 3055 1015
rect 2895 700 2925 800
rect 3025 700 3055 800
rect 2895 465 3055 700
rect 2895 365 2925 465
rect 3025 365 3055 465
rect 2895 140 3055 365
rect 2895 40 2925 140
rect 3025 40 3055 140
rect 2895 15 3055 40
rect 3200 1715 3360 1785
rect 3200 1615 3230 1715
rect 3330 1615 3360 1715
rect 3200 1430 3360 1615
rect 3200 1330 3230 1430
rect 3330 1330 3360 1430
rect 3200 1115 3360 1330
rect 3200 1015 3230 1115
rect 3330 1015 3360 1115
rect 3200 800 3360 1015
rect 3200 700 3230 800
rect 3330 700 3360 800
rect 3200 465 3360 700
rect 3200 365 3230 465
rect 3330 365 3360 465
rect 3200 140 3360 365
rect 3200 40 3230 140
rect 3330 40 3360 140
rect 3200 15 3360 40
rect 3570 1715 3730 1785
rect 3570 1615 3600 1715
rect 3700 1615 3730 1715
rect 3570 1430 3730 1615
rect 3570 1330 3600 1430
rect 3700 1330 3730 1430
rect 3570 1115 3730 1330
rect 3570 1015 3600 1115
rect 3700 1015 3730 1115
rect 3570 800 3730 1015
rect 3570 700 3600 800
rect 3700 700 3730 800
rect 3570 465 3730 700
rect 3570 365 3600 465
rect 3700 365 3730 465
rect 3570 140 3730 365
rect 3875 1715 4035 1785
rect 3875 1615 3905 1715
rect 4005 1615 4035 1715
rect 3875 1430 4035 1615
rect 3875 1330 3905 1430
rect 4005 1330 4035 1430
rect 3875 1115 4035 1330
rect 3875 1015 3905 1115
rect 4005 1015 4035 1115
rect 3875 800 4035 1015
rect 3875 700 3905 800
rect 4005 700 4035 800
rect 3875 465 4035 700
rect 3875 365 3905 465
rect 4005 365 4035 465
rect 3875 140 4035 365
rect 3570 40 3600 140
rect 3700 40 3905 140
rect 4005 40 4035 140
rect 3570 15 3730 40
rect 3875 15 4035 40
rect 4245 1715 4405 1785
rect 4245 1615 4275 1715
rect 4375 1615 4405 1715
rect 4245 1430 4405 1615
rect 4245 1330 4275 1430
rect 4375 1330 4405 1430
rect 4245 1115 4405 1330
rect 4245 1015 4275 1115
rect 4375 1015 4405 1115
rect 4245 800 4405 1015
rect 4245 700 4275 800
rect 4375 700 4405 800
rect 4245 465 4405 700
rect 4245 365 4275 465
rect 4375 365 4405 465
rect 4245 140 4405 365
rect 4245 40 4275 140
rect 4375 40 4405 140
rect 4245 15 4405 40
rect 40 -35 160 -25
rect 40 -135 50 -35
rect 150 -65 160 -35
rect 250 -65 320 15
rect 705 -35 825 -25
rect 705 -65 715 -35
rect 150 -115 715 -65
rect 150 -135 160 -115
rect 40 -145 160 -135
rect 705 -135 715 -115
rect 815 -135 825 -35
rect 705 -145 825 -135
rect 920 -180 970 15
rect 1380 -35 1500 -25
rect 1380 -135 1390 -35
rect 1490 -135 1500 -35
rect 1380 -145 1500 -135
rect 2055 -35 2175 -25
rect 2055 -135 2065 -35
rect 2165 -135 2175 -35
rect 2055 -145 2175 -135
rect 2730 -35 2850 -25
rect 2730 -135 2740 -35
rect 2840 -135 2850 -35
rect 2730 -145 2850 -135
rect 3405 -35 3525 -25
rect 3405 -135 3415 -35
rect 3515 -135 3525 -35
rect 3405 -145 3525 -135
rect 4080 -35 4200 -25
rect 4080 -135 4090 -35
rect 4190 -135 4200 -35
rect 4080 -145 4200 -135
rect 920 -230 1280 -180
rect 40 -385 160 -375
rect 40 -485 50 -385
rect 150 -410 160 -385
rect 705 -385 825 -375
rect 705 -410 715 -385
rect 150 -460 715 -410
rect 150 -485 160 -460
rect 40 -495 160 -485
rect 705 -485 715 -460
rect 815 -485 825 -385
rect 705 -495 825 -485
rect 1230 -410 1280 -230
rect 2095 -255 2145 -145
rect 3415 -180 3515 -145
rect 4335 -210 4385 15
rect 4300 -220 4420 -210
rect 2095 -305 2325 -255
rect 1380 -385 1500 -375
rect 1380 -410 1390 -385
rect 1230 -460 1390 -410
rect 1230 -535 1280 -460
rect 1380 -485 1390 -460
rect 1490 -485 1500 -385
rect 1380 -495 1500 -485
rect 2055 -385 2175 -375
rect 2055 -485 2065 -385
rect 2165 -485 2175 -385
rect 2055 -495 2175 -485
rect 2275 -535 2325 -305
rect 4300 -320 4310 -220
rect 4410 -320 4420 -220
rect 4300 -330 4420 -320
rect 3415 -375 3515 -340
rect 2730 -385 2850 -375
rect 2730 -485 2740 -385
rect 2840 -485 2850 -385
rect 2730 -495 2850 -485
rect 3405 -385 3525 -375
rect 3405 -485 3415 -385
rect 3515 -485 3525 -385
rect 3405 -495 3525 -485
rect 4080 -385 4200 -375
rect 4080 -485 4090 -385
rect 4190 -485 4200 -385
rect 4080 -495 4200 -485
rect 4335 -535 4385 -330
rect -170 -600 -10 -535
rect -170 -700 -140 -600
rect -40 -700 -10 -600
rect -170 -810 -10 -700
rect -170 -910 -140 -810
rect -40 -910 -10 -810
rect -170 -1020 -10 -910
rect -170 -1120 -140 -1020
rect -40 -1120 -10 -1020
rect -170 -1230 -10 -1120
rect -170 -1330 -140 -1230
rect -40 -1330 -10 -1230
rect -170 -1405 -10 -1330
rect 200 -600 360 -535
rect 200 -700 230 -600
rect 330 -700 360 -600
rect 200 -810 360 -700
rect 200 -910 230 -810
rect 330 -910 360 -810
rect 200 -1020 360 -910
rect 200 -1120 230 -1020
rect 330 -1120 360 -1020
rect 200 -1230 360 -1120
rect 200 -1330 230 -1230
rect 330 -1330 360 -1230
rect 200 -1405 360 -1330
rect 500 -600 660 -535
rect 500 -700 530 -600
rect 630 -700 660 -600
rect 500 -810 660 -700
rect 500 -910 530 -810
rect 630 -910 660 -810
rect 500 -1020 660 -910
rect 500 -1120 530 -1020
rect 630 -1120 660 -1020
rect 500 -1230 660 -1120
rect 500 -1330 530 -1230
rect 630 -1330 660 -1230
rect 500 -1405 660 -1330
rect 870 -600 1030 -535
rect 870 -700 900 -600
rect 1000 -700 1030 -600
rect 870 -810 1030 -700
rect 870 -910 900 -810
rect 1000 -910 1030 -810
rect 870 -1020 1030 -910
rect 870 -1120 900 -1020
rect 1000 -1120 1030 -1020
rect 870 -1230 1030 -1120
rect 870 -1330 900 -1230
rect 1000 -1330 1030 -1230
rect 870 -1405 1030 -1330
rect 1175 -600 1335 -535
rect 1175 -700 1205 -600
rect 1305 -700 1335 -600
rect 1175 -810 1335 -700
rect 1175 -910 1205 -810
rect 1305 -910 1335 -810
rect 1175 -1020 1335 -910
rect 1175 -1120 1205 -1020
rect 1305 -1120 1335 -1020
rect 1175 -1230 1335 -1120
rect 1175 -1330 1205 -1230
rect 1305 -1330 1335 -1230
rect 1175 -1405 1335 -1330
rect 1545 -600 1705 -535
rect 1545 -700 1575 -600
rect 1675 -700 1705 -600
rect 1545 -810 1705 -700
rect 1545 -910 1575 -810
rect 1675 -910 1705 -810
rect 1545 -1020 1705 -910
rect 1545 -1120 1575 -1020
rect 1675 -1120 1705 -1020
rect 1545 -1230 1705 -1120
rect 1545 -1330 1575 -1230
rect 1675 -1330 1705 -1230
rect 1545 -1405 1705 -1330
rect 1850 -600 2010 -535
rect 1850 -700 1880 -600
rect 1980 -700 2010 -600
rect 1850 -810 2010 -700
rect 1850 -910 1880 -810
rect 1980 -910 2010 -810
rect 1850 -1020 2010 -910
rect 1850 -1120 1880 -1020
rect 1980 -1120 2010 -1020
rect 1850 -1230 2010 -1120
rect 1850 -1330 1880 -1230
rect 1980 -1330 2010 -1230
rect 1850 -1405 2010 -1330
rect 2220 -600 2380 -535
rect 2220 -700 2250 -600
rect 2350 -700 2380 -600
rect 2220 -810 2380 -700
rect 2220 -910 2250 -810
rect 2350 -910 2380 -810
rect 2220 -1020 2380 -910
rect 2220 -1120 2250 -1020
rect 2350 -1120 2380 -1020
rect 2220 -1230 2380 -1120
rect 2220 -1330 2250 -1230
rect 2350 -1330 2380 -1230
rect 2220 -1405 2380 -1330
rect 2525 -600 2685 -535
rect 2525 -700 2555 -600
rect 2655 -700 2685 -600
rect 2525 -810 2685 -700
rect 2525 -910 2555 -810
rect 2655 -910 2685 -810
rect 2525 -1020 2685 -910
rect 2525 -1120 2555 -1020
rect 2655 -1120 2685 -1020
rect 2525 -1230 2685 -1120
rect 2525 -1330 2555 -1230
rect 2655 -1330 2685 -1230
rect 2525 -1405 2685 -1330
rect 2895 -600 3055 -535
rect 2895 -700 2925 -600
rect 3025 -700 3055 -600
rect 2895 -810 3055 -700
rect 2895 -910 2925 -810
rect 3025 -910 3055 -810
rect 2895 -1020 3055 -910
rect 2895 -1120 2925 -1020
rect 3025 -1120 3055 -1020
rect 2895 -1230 3055 -1120
rect 2895 -1330 2925 -1230
rect 3025 -1305 3055 -1230
rect 3200 -600 3360 -535
rect 3200 -700 3230 -600
rect 3330 -700 3360 -600
rect 3200 -810 3360 -700
rect 3200 -910 3230 -810
rect 3330 -910 3360 -810
rect 3200 -1020 3360 -910
rect 3200 -1120 3230 -1020
rect 3330 -1120 3360 -1020
rect 3200 -1230 3360 -1120
rect 3200 -1305 3230 -1230
rect 3025 -1330 3230 -1305
rect 3330 -1330 3360 -1230
rect 2895 -1405 3360 -1330
rect 3570 -600 3730 -535
rect 3570 -700 3600 -600
rect 3700 -605 3730 -600
rect 3875 -600 4035 -535
rect 3875 -605 3905 -600
rect 3700 -700 3905 -605
rect 4005 -700 4035 -600
rect 3570 -705 4035 -700
rect 3570 -810 3730 -705
rect 3570 -910 3600 -810
rect 3700 -910 3730 -810
rect 3570 -1020 3730 -910
rect 3570 -1120 3600 -1020
rect 3700 -1120 3730 -1020
rect 3570 -1230 3730 -1120
rect 3570 -1330 3600 -1230
rect 3700 -1330 3730 -1230
rect 3570 -1405 3730 -1330
rect 3875 -810 4035 -705
rect 3875 -910 3905 -810
rect 4005 -910 4035 -810
rect 3875 -1020 4035 -910
rect 3875 -1120 3905 -1020
rect 4005 -1120 4035 -1020
rect 3875 -1230 4035 -1120
rect 3875 -1330 3905 -1230
rect 4005 -1330 4035 -1230
rect 3875 -1405 4035 -1330
rect 4245 -600 4405 -535
rect 4245 -700 4275 -600
rect 4375 -700 4405 -600
rect 4245 -810 4405 -700
rect 4245 -910 4275 -810
rect 4375 -910 4405 -810
rect 4245 -1020 4405 -910
rect 4245 -1120 4275 -1020
rect 4375 -1120 4405 -1020
rect 4245 -1230 4405 -1120
rect 4245 -1330 4275 -1230
rect 4375 -1330 4405 -1230
rect 4245 -1405 4405 -1330
rect -155 -1540 -20 -1405
rect -155 -1650 -145 -1540
rect -30 -1650 -20 -1540
rect -155 -1660 -20 -1650
rect 515 -1540 650 -1405
rect 515 -1650 525 -1540
rect 640 -1650 650 -1540
rect 515 -1660 650 -1650
rect 2050 -1540 2185 -1530
rect 2050 -1650 2060 -1540
rect 2175 -1650 2185 -1540
rect 2050 -1660 2185 -1650
rect 2910 -1540 3045 -1405
rect 2910 -1650 2920 -1540
rect 3035 -1650 3045 -1540
rect 3405 -1460 3525 -1450
rect 3405 -1560 3415 -1460
rect 3515 -1560 3525 -1460
rect 3405 -1570 3525 -1560
rect 2910 -1660 3045 -1650
<< viali >>
rect -145 1890 -30 2000
rect 525 1890 640 2000
rect 2060 1885 2175 1995
rect 2915 1890 3030 2000
rect 230 40 330 140
rect 1205 40 1305 140
rect 1575 700 1675 800
rect 1880 700 1980 800
rect 2250 365 2350 465
rect 2250 45 2350 145
rect 2555 700 2655 800
rect 2925 365 3025 465
rect 1390 -135 1490 -35
rect 2740 -135 2840 -35
rect 4090 -135 4190 -35
rect 1390 -485 1490 -385
rect 2065 -485 2165 -385
rect 4310 -320 4410 -220
rect 2740 -485 2840 -385
rect 4090 -485 4190 -385
rect 230 -700 330 -600
rect 900 -700 1000 -600
rect 1575 -700 1675 -600
rect 1880 -700 1980 -600
rect 2250 -910 2350 -810
rect 2555 -700 2655 -600
rect 2925 -910 3025 -810
rect -145 -1650 -30 -1540
rect 525 -1650 640 -1540
rect 2060 -1650 2175 -1540
rect 2920 -1650 3035 -1540
<< metal1 >>
rect -155 2000 -20 2010
rect -155 1890 -145 2000
rect -30 1890 -20 2000
rect -155 1880 -20 1890
rect 515 2000 650 2010
rect 515 1890 525 2000
rect 640 1890 650 2000
rect 515 1880 650 1890
rect 2050 1995 2185 2005
rect 2050 1885 2060 1995
rect 2175 1885 2185 1995
rect 2050 1880 2185 1885
rect 2905 2000 3040 2010
rect 2905 1890 2915 2000
rect 3030 1890 3040 2000
rect 2905 1880 3040 1890
rect 1565 800 2665 810
rect 1565 700 1575 800
rect 1675 700 1880 800
rect 1980 700 2555 800
rect 2655 700 2665 800
rect 1565 690 2665 700
rect 2240 465 3035 475
rect 2240 365 2250 465
rect 2350 365 2925 465
rect 3025 365 3035 465
rect 2240 355 3035 365
rect 220 140 340 150
rect 220 40 230 140
rect 330 40 340 140
rect 220 30 340 40
rect 1195 140 1315 150
rect 1195 40 1205 140
rect 1305 40 1315 140
rect 1195 30 1315 40
rect 2240 145 2360 155
rect 2240 45 2250 145
rect 2350 45 2360 145
rect 2240 35 2360 45
rect 260 -590 310 30
rect 1230 -95 1280 30
rect 1380 -35 1500 -25
rect 1380 -95 1390 -35
rect 1230 -135 1390 -95
rect 1490 -135 1500 -35
rect 1230 -145 1500 -135
rect 1230 -330 1280 -145
rect 2275 -215 2325 35
rect 920 -380 1280 -330
rect 2095 -265 2325 -215
rect 2730 -35 2850 -25
rect 2730 -135 2740 -35
rect 2840 -135 2850 -35
rect 2730 -210 2850 -135
rect 4080 -35 4200 -25
rect 4080 -135 4090 -35
rect 4190 -135 4200 -35
rect 4080 -145 4200 -135
rect 2730 -220 4420 -210
rect 2095 -375 2145 -265
rect 2730 -320 4310 -220
rect 4410 -320 4420 -220
rect 2730 -330 4420 -320
rect 920 -590 970 -380
rect 1380 -385 1500 -375
rect 1380 -485 1390 -385
rect 1490 -485 1500 -385
rect 1380 -495 1500 -485
rect 2055 -385 2175 -375
rect 2055 -485 2065 -385
rect 2165 -485 2175 -385
rect 2055 -490 2175 -485
rect 2730 -385 2850 -330
rect 2730 -485 2740 -385
rect 2840 -485 2850 -385
rect 2730 -495 2850 -485
rect 4080 -385 4200 -375
rect 4080 -485 4090 -385
rect 4190 -485 4200 -385
rect 4080 -495 4200 -485
rect 220 -600 340 -590
rect 220 -700 230 -600
rect 330 -700 340 -600
rect 220 -710 340 -700
rect 890 -600 1010 -590
rect 890 -700 900 -600
rect 1000 -700 1010 -600
rect 890 -710 1010 -700
rect 1565 -600 2665 -590
rect 1565 -700 1575 -600
rect 1675 -700 1880 -600
rect 1980 -700 2555 -600
rect 2655 -700 2665 -600
rect 1565 -710 2665 -700
rect 2240 -810 3035 -800
rect 2240 -910 2250 -810
rect 2350 -910 2925 -810
rect 3025 -910 3035 -810
rect 2240 -920 3035 -910
rect -155 -1540 -20 -1530
rect -155 -1650 -145 -1540
rect -30 -1650 -20 -1540
rect -155 -1660 -20 -1650
rect 515 -1540 650 -1530
rect 515 -1650 525 -1540
rect 640 -1650 650 -1540
rect 515 -1660 650 -1650
rect 2050 -1540 2185 -1530
rect 2050 -1650 2060 -1540
rect 2175 -1650 2185 -1540
rect 2050 -1660 2185 -1650
rect 2910 -1540 3045 -1530
rect 2910 -1650 2920 -1540
rect 3035 -1650 3045 -1540
rect 2910 -1660 3045 -1650
<< via1 >>
rect -145 1890 -30 2000
rect 525 1890 640 2000
rect 2060 1885 2175 1995
rect 2915 1890 3030 2000
rect 1390 -135 1490 -35
rect 4090 -135 4190 -35
rect 1390 -485 1490 -385
rect 4090 -485 4190 -385
rect -145 -1650 -30 -1540
rect 525 -1650 640 -1540
rect 2060 -1650 2175 -1540
rect 2920 -1650 3035 -1540
<< metal2 >>
rect -155 2000 -20 2010
rect -155 1890 -145 2000
rect -30 1890 -20 2000
rect -155 1880 -20 1890
rect 515 2000 650 2010
rect 515 1890 525 2000
rect 640 1890 650 2000
rect 515 1880 650 1890
rect 2050 1995 2185 2005
rect 2050 1885 2060 1995
rect 2175 1885 2185 1995
rect 2050 1880 2185 1885
rect 2905 2000 3040 2010
rect 2905 1890 2915 2000
rect 3030 1890 3040 2000
rect 2905 1880 3040 1890
rect 1380 -35 1500 -25
rect 1380 -135 1390 -35
rect 1490 -135 1500 -35
rect 1380 -145 1500 -135
rect 4080 -35 4200 -25
rect 4080 -135 4090 -35
rect 4190 -135 4200 -35
rect 4080 -145 4200 -135
rect 1380 -385 1500 -375
rect 4080 -385 4200 -375
rect 1380 -485 1390 -385
rect 1490 -485 4090 -385
rect 4190 -485 4200 -385
rect 1380 -495 1500 -485
rect 4080 -495 4200 -485
rect -155 -1540 -20 -1530
rect -155 -1650 -145 -1540
rect -30 -1650 -20 -1540
rect -155 -1660 -20 -1650
rect 515 -1540 650 -1530
rect 515 -1650 525 -1540
rect 640 -1650 650 -1540
rect 515 -1660 650 -1650
rect 2050 -1540 2185 -1530
rect 2050 -1650 2060 -1540
rect 2175 -1650 2185 -1540
rect 2050 -1660 2185 -1650
rect 2910 -1540 3045 -1530
rect 2910 -1650 2920 -1540
rect 3035 -1650 3045 -1540
rect 2910 -1660 3045 -1650
<< via2 >>
rect -145 1890 -30 2000
rect 525 1890 640 2000
rect 2060 1885 2175 1995
rect 2915 1890 3030 2000
rect 1390 -135 1490 -35
rect 4090 -135 4190 -35
rect -145 -1650 -30 -1540
rect 525 -1650 640 -1540
rect 2060 -1650 2175 -1540
rect 2920 -1650 3035 -1540
<< metal3 >>
rect -155 2000 -20 2010
rect -155 1890 -145 2000
rect -30 1890 -20 2000
rect -155 1880 -20 1890
rect 515 2000 650 2010
rect 515 1890 525 2000
rect 640 1890 650 2000
rect 515 1880 650 1890
rect 2050 1995 2185 2005
rect 2050 1885 2060 1995
rect 2175 1885 2185 1995
rect 2050 1880 2185 1885
rect 2905 2000 3040 2010
rect 2905 1890 2915 2000
rect 3030 1890 3040 2000
rect 2905 1880 3040 1890
rect 1380 -35 1500 -25
rect 4080 -35 4200 -25
rect 1380 -135 1390 -35
rect 1490 -135 4090 -35
rect 4190 -135 4200 -35
rect 1380 -145 1500 -135
rect 4080 -145 4200 -135
rect -155 -1540 -20 -1530
rect -155 -1650 -145 -1540
rect -30 -1650 -20 -1540
rect -155 -1660 -20 -1650
rect 515 -1540 650 -1530
rect 515 -1650 525 -1540
rect 640 -1650 650 -1540
rect 515 -1660 650 -1650
rect 2050 -1540 2185 -1530
rect 2050 -1650 2060 -1540
rect 2175 -1650 2185 -1540
rect 2050 -1660 2185 -1650
rect 2910 -1540 3045 -1530
rect 2910 -1650 2920 -1540
rect 3035 -1650 3045 -1540
rect 2910 -1660 3045 -1650
<< via3 >>
rect -145 1890 -30 2000
rect 525 1890 640 2000
rect 2060 1885 2175 1995
rect 2915 1890 3030 2000
rect -145 -1650 -30 -1540
rect 525 -1650 640 -1540
rect 2060 -1650 2175 -1540
rect 2920 -1650 3035 -1540
<< metal4 >>
rect -245 2000 4500 2030
rect -245 1890 -145 2000
rect -30 1890 525 2000
rect 640 1995 2915 2000
rect 640 1890 2060 1995
rect -245 1885 2060 1890
rect 2175 1890 2915 1995
rect 3030 1890 4500 2000
rect 2175 1885 4500 1890
rect -245 1860 4500 1885
rect -245 -1540 4495 -1475
rect -245 -1650 -145 -1540
rect -30 -1650 525 -1540
rect 640 -1650 2060 -1540
rect 2175 -1650 2920 -1540
rect 3035 -1650 4495 -1540
rect -245 -1715 4495 -1650
<< labels >>
rlabel locali 430 -435 430 -435 1 vbias
rlabel locali 2115 1995 2115 1995 1 vdd!
rlabel locali 2140 -1650 2140 -1650 1 gnd!
rlabel locali 4360 -155 4360 -155 1 out
rlabel locali 3465 -360 3465 -360 1 down
rlabel locali 3465 -160 3465 -160 1 upbar
<< end >>
