magic
tech sky130A
magscale 1 2
timestamp 1640901950
<< error_s >>
rect 764 1710 855 2110
rect 7081 1710 7154 2110
rect 1616 -3178 1796 -2353
rect 1616 -6718 1796 -5278
rect 1616 -10288 1796 -8848
<< psubdiff >>
rect 8630 150 8890 180
rect 8630 -50 8660 150
rect 8860 -50 8890 150
rect 8630 -80 8890 -50
rect 8630 -510 8890 -480
rect 8630 -710 8660 -510
rect 8860 -710 8890 -510
rect 8630 -740 8890 -710
rect 8630 -1170 8890 -1140
rect 8630 -1370 8660 -1170
rect 8860 -1370 8890 -1170
rect 8630 -1400 8890 -1370
rect 8630 -1830 8890 -1800
rect 8630 -2030 8660 -1830
rect 8860 -2030 8890 -1830
rect 8630 -2060 8890 -2030
rect 8630 -2490 8890 -2460
rect 8630 -2690 8660 -2490
rect 8860 -2690 8890 -2490
rect 8630 -2720 8890 -2690
rect 8630 -3150 8890 -3120
rect 8630 -3350 8660 -3150
rect 8860 -3350 8890 -3150
rect 8630 -3380 8890 -3350
rect 8630 -3810 8890 -3780
rect 8630 -4010 8660 -3810
rect 8860 -4010 8890 -3810
rect 8630 -4040 8890 -4010
rect 8630 -4470 8890 -4440
rect 8630 -4670 8660 -4470
rect 8860 -4670 8890 -4470
rect 8630 -4700 8890 -4670
rect 8630 -5130 8890 -5100
rect 8630 -5330 8660 -5130
rect 8860 -5330 8890 -5130
rect 8630 -5360 8890 -5330
rect 8630 -5790 8890 -5760
rect 8630 -5990 8660 -5790
rect 8860 -5990 8890 -5790
rect 8630 -6020 8890 -5990
rect 8630 -6450 8890 -6420
rect 8630 -6650 8660 -6450
rect 8860 -6650 8890 -6450
rect 8630 -6680 8890 -6650
rect 8630 -7110 8890 -7080
rect 8630 -7310 8660 -7110
rect 8860 -7310 8890 -7110
rect 8630 -7340 8890 -7310
rect 8630 -7770 8890 -7740
rect 8630 -7970 8660 -7770
rect 8860 -7970 8890 -7770
rect 8630 -8000 8890 -7970
rect 8630 -8430 8890 -8400
rect 8630 -8630 8660 -8430
rect 8860 -8630 8890 -8430
rect 8630 -8660 8890 -8630
rect 8630 -9090 8890 -9060
rect 8630 -9290 8660 -9090
rect 8860 -9290 8890 -9090
rect 8630 -9320 8890 -9290
rect 8630 -9750 8890 -9720
rect 8630 -9950 8660 -9750
rect 8860 -9950 8890 -9750
rect 8630 -9980 8890 -9950
rect 7790 -10410 8050 -10380
rect 7790 -10610 7820 -10410
rect 8020 -10610 8050 -10410
rect 7790 -10640 8050 -10610
rect 8630 -10410 8890 -10380
rect 8630 -10610 8660 -10410
rect 8860 -10610 8890 -10410
rect 8630 -10640 8890 -10610
<< psubdiffcont >>
rect 8660 -50 8860 150
rect 8660 -710 8860 -510
rect 8660 -1370 8860 -1170
rect 8660 -2030 8860 -1830
rect 8660 -2690 8860 -2490
rect 8660 -3350 8860 -3150
rect 8660 -4010 8860 -3810
rect 8660 -4670 8860 -4470
rect 8660 -5330 8860 -5130
rect 8660 -5990 8860 -5790
rect 8660 -6650 8860 -6450
rect 8660 -7310 8860 -7110
rect 8660 -7970 8860 -7770
rect 8660 -8630 8860 -8430
rect 8660 -9290 8860 -9090
rect 8660 -9950 8860 -9750
rect 7820 -10610 8020 -10410
rect 8660 -10610 8860 -10410
<< locali >>
rect 7440 1500 7620 1520
rect 1330 1480 1470 1500
rect 1330 1460 1350 1480
rect 1010 1400 1350 1460
rect 1330 1380 1350 1400
rect 1450 1380 1470 1480
rect 4420 1470 4560 1490
rect 4420 1450 4440 1470
rect 4080 1390 4440 1450
rect 1330 1360 1470 1380
rect 4420 1370 4440 1390
rect 4540 1370 4560 1470
rect 7440 1460 7460 1500
rect 7140 1400 7460 1460
rect 4420 1350 4560 1370
rect 7440 1360 7460 1400
rect 7600 1360 7620 1500
rect 7440 1340 7620 1360
rect 8640 150 8880 170
rect 8640 -50 8660 150
rect 8860 -50 8880 150
rect 8640 -70 8880 -50
rect 8640 -510 8880 -490
rect 8640 -710 8660 -510
rect 8860 -710 8880 -510
rect 8640 -730 8880 -710
rect 8640 -1170 8880 -1150
rect 8640 -1370 8660 -1170
rect 8860 -1370 8880 -1170
rect 8640 -1390 8880 -1370
rect 1916 -1680 2286 -1610
rect 2924 -1680 3264 -1610
rect 3872 -1680 4242 -1610
rect 4852 -1680 5212 -1610
rect 5834 -1680 6194 -1610
rect 6856 -1680 7386 -1610
rect 2216 -5150 2286 -1680
rect 3194 -5150 3264 -1680
rect 4172 -5150 4242 -1680
rect 5142 -5150 5212 -1680
rect 6124 -5150 6194 -1680
rect 7316 -5150 7386 -1680
rect 8640 -1830 8880 -1810
rect 8640 -2030 8660 -1830
rect 8860 -2030 8880 -1830
rect 8640 -2050 8880 -2030
rect 8640 -2490 8880 -2470
rect 8640 -2690 8660 -2490
rect 8860 -2690 8880 -2490
rect 8640 -2710 8880 -2690
rect 8640 -3150 8880 -3130
rect 8640 -3350 8660 -3150
rect 8860 -3350 8880 -3150
rect 8640 -3370 8880 -3350
rect 8640 -3810 8880 -3790
rect 8640 -4010 8660 -3810
rect 8860 -4010 8880 -3810
rect 8640 -4030 8880 -4010
rect 8640 -4470 8880 -4450
rect 8640 -4670 8660 -4470
rect 8860 -4670 8880 -4470
rect 8640 -4690 8880 -4670
rect 1916 -5220 2286 -5150
rect 2924 -5220 3264 -5150
rect 3872 -5220 4242 -5150
rect 4852 -5220 5212 -5150
rect 5834 -5220 6194 -5150
rect 6856 -5220 7386 -5150
rect 2216 -8720 2286 -5220
rect 3194 -8720 3264 -5220
rect 4172 -8720 4242 -5220
rect 5142 -8720 5212 -5220
rect 6124 -8720 6194 -5220
rect 7316 -8720 7386 -5220
rect 8640 -5130 8880 -5110
rect 8640 -5330 8660 -5130
rect 8860 -5330 8880 -5130
rect 8640 -5350 8880 -5330
rect 8640 -5790 8880 -5770
rect 8640 -5990 8660 -5790
rect 8860 -5990 8880 -5790
rect 8640 -6010 8880 -5990
rect 8640 -6450 8880 -6430
rect 8640 -6650 8660 -6450
rect 8860 -6650 8880 -6450
rect 8640 -6670 8880 -6650
rect 8640 -7110 8880 -7090
rect 8640 -7310 8660 -7110
rect 8860 -7310 8880 -7110
rect 8640 -7330 8880 -7310
rect 8640 -7770 8880 -7750
rect 8640 -7970 8660 -7770
rect 8860 -7970 8880 -7770
rect 8640 -7990 8880 -7970
rect 8640 -8430 8880 -8410
rect 8640 -8630 8660 -8430
rect 8860 -8630 8880 -8430
rect 8640 -8650 8880 -8630
rect 1916 -8790 2286 -8720
rect 2924 -8790 3264 -8720
rect 3872 -8790 4242 -8720
rect 4852 -8790 5212 -8720
rect 5834 -8790 6194 -8720
rect 6856 -8790 7386 -8720
rect 8640 -9090 8880 -9070
rect 8640 -9290 8660 -9090
rect 8860 -9290 8880 -9090
rect 8640 -9310 8880 -9290
rect 8640 -9750 8880 -9730
rect 8640 -9950 8660 -9750
rect 8860 -9950 8880 -9750
rect 8640 -9970 8880 -9950
rect 7800 -10410 8040 -10390
rect 7800 -10610 7820 -10410
rect 8020 -10610 8040 -10410
rect 7800 -10630 8040 -10610
rect 8640 -10410 8880 -10390
rect 8640 -10610 8660 -10410
rect 8860 -10610 8880 -10410
rect 8640 -10630 8880 -10610
<< viali >>
rect 1350 1380 1450 1480
rect 4440 1370 4540 1470
rect 7460 1360 7600 1500
rect 8660 -50 8860 150
rect 8660 -710 8860 -510
rect 8660 -1370 8860 -1170
rect 8660 -2030 8860 -1830
rect 8660 -2690 8860 -2490
rect 8660 -3350 8860 -3150
rect 8660 -4010 8860 -3810
rect 8660 -4670 8860 -4470
rect 8660 -5330 8860 -5130
rect 8660 -5990 8860 -5790
rect 8660 -6650 8860 -6450
rect 8660 -7310 8860 -7110
rect 8660 -7970 8860 -7770
rect 8660 -8630 8860 -8430
rect 8660 -9290 8860 -9090
rect 8660 -9950 8860 -9750
rect 7820 -10610 8020 -10410
rect 8660 -10610 8860 -10410
<< metal1 >>
rect 7440 1500 7620 1520
rect 1330 1480 1470 1500
rect 1330 1380 1350 1480
rect 1450 1380 1470 1480
rect 1330 1360 1470 1380
rect 4420 1470 4560 1490
rect 4420 1370 4440 1470
rect 4540 1370 4560 1470
rect 4420 1350 4560 1370
rect 7440 1360 7460 1500
rect 7600 1360 7620 1500
rect 7440 1340 7620 1360
rect 8650 860 8870 870
rect 8650 850 8660 860
rect 7180 670 8660 850
rect 8650 660 8660 670
rect 8860 660 8870 860
rect 8650 650 8870 660
rect 8640 150 8880 170
rect 8640 -50 8660 150
rect 8860 -50 8880 150
rect 8640 -70 8880 -50
rect 8640 -510 8880 -490
rect 8640 -710 8660 -510
rect 8860 -710 8880 -510
rect 8640 -730 8880 -710
rect 8640 -1170 8880 -1150
rect 8640 -1370 8660 -1170
rect 8860 -1370 8880 -1170
rect 8640 -1390 8880 -1370
rect 8640 -1830 8880 -1810
rect 8640 -2030 8660 -1830
rect 8860 -2030 8880 -1830
rect 8640 -2050 8880 -2030
rect 8640 -2490 8880 -2470
rect 8640 -2690 8660 -2490
rect 8860 -2690 8880 -2490
rect 8640 -2710 8880 -2690
rect 8640 -3150 8880 -3130
rect 8640 -3350 8660 -3150
rect 8860 -3350 8880 -3150
rect 8640 -3370 8880 -3350
rect 8640 -3810 8880 -3790
rect 8640 -4010 8660 -3810
rect 8860 -4010 8880 -3810
rect 8640 -4030 8880 -4010
rect 8640 -4470 8880 -4450
rect 8640 -4670 8660 -4470
rect 8860 -4670 8880 -4470
rect 8640 -4690 8880 -4670
rect 8640 -5130 8880 -5110
rect 8640 -5330 8660 -5130
rect 8860 -5330 8880 -5130
rect 8640 -5350 8880 -5330
rect 8640 -5790 8880 -5770
rect 8640 -5990 8660 -5790
rect 8860 -5990 8880 -5790
rect 8640 -6010 8880 -5990
rect 8640 -6450 8880 -6430
rect 8640 -6650 8660 -6450
rect 8860 -6650 8880 -6450
rect 8640 -6670 8880 -6650
rect 8640 -7110 8880 -7090
rect 8640 -7310 8660 -7110
rect 8860 -7310 8880 -7110
rect 8640 -7330 8880 -7310
rect 8640 -7770 8880 -7750
rect 8640 -7970 8660 -7770
rect 8860 -7970 8880 -7770
rect 8640 -7990 8880 -7970
rect 8640 -8430 8880 -8410
rect 8640 -8630 8660 -8430
rect 8860 -8630 8880 -8430
rect 8640 -8650 8880 -8630
rect 8640 -9090 8880 -9070
rect 8640 -9290 8660 -9090
rect 8860 -9290 8880 -9090
rect 8640 -9310 8880 -9290
rect 8640 -9750 8880 -9730
rect 8640 -9950 8660 -9750
rect 8860 -9950 8880 -9750
rect 8640 -9970 8880 -9950
rect 7800 -10410 8040 -10390
rect 7800 -10610 7820 -10410
rect 8020 -10610 8040 -10410
rect 7800 -10630 8040 -10610
rect 8640 -10410 8880 -10390
rect 8640 -10610 8660 -10410
rect 8860 -10610 8880 -10410
rect 8640 -10630 8880 -10610
<< via1 >>
rect 1350 1380 1450 1480
rect 4440 1370 4540 1470
rect 7460 1360 7600 1500
rect 8660 660 8860 860
rect 8660 -50 8860 150
rect 8660 -710 8860 -510
rect 8660 -1370 8860 -1170
rect 8660 -2030 8860 -1830
rect 8660 -2690 8860 -2490
rect 8660 -3350 8860 -3150
rect 8660 -4010 8860 -3810
rect 8660 -4670 8860 -4470
rect 8660 -5330 8860 -5130
rect 8660 -5990 8860 -5790
rect 8660 -6650 8860 -6450
rect 8660 -7310 8860 -7110
rect 8660 -7970 8860 -7770
rect 8660 -8630 8860 -8430
rect 8660 -9290 8860 -9090
rect 8660 -9950 8860 -9750
rect 7820 -10610 8020 -10410
rect 8660 -10610 8860 -10410
<< metal2 >>
rect 7420 1500 8240 1550
rect 1330 1480 1470 1500
rect 1330 1380 1350 1480
rect 1450 1380 1470 1480
rect 1330 1360 1470 1380
rect 4420 1470 4560 1490
rect 4420 1370 4440 1470
rect 4540 1370 4560 1470
rect 4420 1350 4560 1370
rect 7420 1360 7460 1500
rect 7600 1360 8240 1500
rect 7420 1310 8240 1360
rect 8000 -7410 8240 1310
rect 8650 860 8870 870
rect 8650 660 8660 860
rect 8860 660 8870 860
rect 8650 650 8870 660
rect 8640 150 8880 170
rect 8640 -50 8660 150
rect 8860 -50 8880 150
rect 8640 -70 8880 -50
rect 8640 -510 8880 -490
rect 8640 -710 8660 -510
rect 8860 -710 8880 -510
rect 8640 -730 8880 -710
rect 8640 -1170 8880 -1150
rect 8640 -1370 8660 -1170
rect 8860 -1370 8880 -1170
rect 8640 -1390 8880 -1370
rect 8640 -1830 8880 -1810
rect 8640 -2030 8660 -1830
rect 8860 -2030 8880 -1830
rect 8640 -2050 8880 -2030
rect 8640 -2490 8880 -2470
rect 8640 -2690 8660 -2490
rect 8860 -2690 8880 -2490
rect 8640 -2710 8880 -2690
rect 8640 -3150 8880 -3130
rect 8640 -3350 8660 -3150
rect 8860 -3350 8880 -3150
rect 8640 -3370 8880 -3350
rect 8640 -3810 8880 -3790
rect 8640 -4010 8660 -3810
rect 8860 -4010 8880 -3810
rect 8640 -4030 8880 -4010
rect 8640 -4470 8880 -4450
rect 8640 -4670 8660 -4470
rect 8860 -4670 8880 -4470
rect 8640 -4690 8880 -4670
rect 8640 -5130 8880 -5110
rect 8640 -5330 8660 -5130
rect 8860 -5330 8880 -5130
rect 8640 -5350 8880 -5330
rect 8640 -5790 8880 -5770
rect 8640 -5990 8660 -5790
rect 8860 -5990 8880 -5790
rect 8640 -6010 8880 -5990
rect 8640 -6450 8880 -6430
rect 8640 -6650 8660 -6450
rect 8860 -6650 8880 -6450
rect 8640 -6670 8880 -6650
rect 8640 -7110 8880 -7090
rect 8640 -7310 8660 -7110
rect 8860 -7310 8880 -7110
rect 8640 -7330 8880 -7310
rect 6916 -7430 8240 -7410
rect 6916 -7630 6936 -7430
rect 7136 -7630 8240 -7430
rect 6916 -7650 8240 -7630
rect 8640 -7770 8880 -7750
rect 8640 -7970 8660 -7770
rect 8860 -7970 8880 -7770
rect 8640 -7990 8880 -7970
rect 8640 -8430 8880 -8410
rect 8640 -8630 8660 -8430
rect 8860 -8630 8880 -8430
rect 8640 -8650 8880 -8630
rect 8640 -9090 8880 -9070
rect 8640 -9290 8660 -9090
rect 8860 -9290 8880 -9090
rect 8640 -9310 8880 -9290
rect 8640 -9750 8880 -9730
rect 8640 -9950 8660 -9750
rect 8860 -9950 8880 -9750
rect 8640 -9970 8880 -9950
rect 7800 -10410 8040 -10390
rect 7800 -10610 7820 -10410
rect 8020 -10610 8040 -10410
rect 7800 -10630 8040 -10610
rect 8640 -10410 8880 -10390
rect 8640 -10610 8660 -10410
rect 8860 -10610 8880 -10410
rect 8640 -10630 8880 -10610
<< via2 >>
rect 1350 1380 1450 1480
rect 4440 1370 4540 1470
rect 8660 660 8860 860
rect 8660 -50 8860 150
rect 8660 -710 8860 -510
rect 8660 -1370 8860 -1170
rect 8660 -2030 8860 -1830
rect 8660 -2690 8860 -2490
rect 8660 -3350 8860 -3150
rect 8660 -4010 8860 -3810
rect 8660 -4670 8860 -4470
rect 8660 -5330 8860 -5130
rect 8660 -5990 8860 -5790
rect 8660 -6650 8860 -6450
rect 8660 -7310 8860 -7110
rect 6936 -7630 7136 -7430
rect 8660 -7970 8860 -7770
rect 8660 -8630 8860 -8430
rect 8660 -9290 8860 -9090
rect 8660 -9950 8860 -9750
rect 7820 -10610 8020 -10410
rect 8660 -10610 8860 -10410
<< metal3 >>
rect 1330 1480 1470 1500
rect 1330 1380 1350 1480
rect 1450 1380 1470 1480
rect 1330 1360 1470 1380
rect 4390 1470 4590 1520
rect 4390 1370 4440 1470
rect 4540 1370 4590 1470
rect 4390 420 4590 1370
rect 8650 860 8870 870
rect 8650 660 8660 860
rect 8860 660 8870 860
rect 8650 650 8870 660
rect 4390 220 7780 420
rect 7580 -3840 7780 220
rect 8640 150 8880 170
rect 8640 -50 8660 150
rect 8860 -50 8880 150
rect 8640 -70 8880 -50
rect 8640 -510 8880 -490
rect 8640 -710 8660 -510
rect 8860 -710 8880 -510
rect 8640 -730 8880 -710
rect 8640 -1170 8880 -1150
rect 8640 -1370 8660 -1170
rect 8860 -1370 8880 -1170
rect 8640 -1390 8880 -1370
rect 8640 -1830 8880 -1810
rect 8640 -2030 8660 -1830
rect 8860 -2030 8880 -1830
rect 8640 -2050 8880 -2030
rect 8640 -2490 8880 -2470
rect 8640 -2690 8660 -2490
rect 8860 -2690 8880 -2490
rect 8640 -2710 8880 -2690
rect 8640 -3150 8880 -3130
rect 8640 -3350 8660 -3150
rect 8860 -3350 8880 -3150
rect 8640 -3370 8880 -3350
rect 6906 -3860 7780 -3840
rect 6906 -4060 6926 -3860
rect 7126 -4060 7780 -3860
rect 8640 -3810 8880 -3790
rect 8640 -4010 8660 -3810
rect 8860 -4010 8880 -3810
rect 8640 -4030 8880 -4010
rect 6906 -4080 7780 -4060
rect 8640 -4470 8880 -4450
rect 8640 -4670 8660 -4470
rect 8860 -4670 8880 -4470
rect 8640 -4690 8880 -4670
rect 8640 -5130 8880 -5110
rect 8640 -5330 8660 -5130
rect 8860 -5330 8880 -5130
rect 8640 -5350 8880 -5330
rect 8640 -5790 8880 -5770
rect 8640 -5990 8660 -5790
rect 8860 -5990 8880 -5790
rect 8640 -6010 8880 -5990
rect 8640 -6450 8880 -6430
rect 8640 -6650 8660 -6450
rect 8860 -6650 8880 -6450
rect 8640 -6670 8880 -6650
rect 8640 -7110 8880 -7090
rect 8640 -7310 8660 -7110
rect 8860 -7310 8880 -7110
rect 8640 -7330 8880 -7310
rect 6916 -7430 7156 -7410
rect 6916 -7630 6936 -7430
rect 7136 -7630 7156 -7430
rect 6916 -7650 7156 -7630
rect 8640 -7770 8880 -7750
rect 8640 -7970 8660 -7770
rect 8860 -7970 8880 -7770
rect 8640 -7990 8880 -7970
rect 8640 -8430 8880 -8410
rect 8640 -8630 8660 -8430
rect 8860 -8630 8880 -8430
rect 8640 -8650 8880 -8630
rect 8640 -9090 8880 -9070
rect 8640 -9290 8660 -9090
rect 8860 -9290 8880 -9090
rect 8640 -9310 8880 -9290
rect 8640 -9750 8880 -9730
rect 8640 -9950 8660 -9750
rect 8860 -9950 8880 -9750
rect 8640 -9970 8880 -9950
rect 7800 -10410 8040 -10390
rect 7800 -10610 7820 -10410
rect 8020 -10610 8040 -10410
rect 7800 -10630 8040 -10610
rect 8640 -10410 8880 -10390
rect 8640 -10610 8660 -10410
rect 8860 -10610 8880 -10410
rect 8640 -10630 8880 -10610
<< via3 >>
rect 1350 1380 1450 1480
rect 8660 660 8860 860
rect 8660 -50 8860 150
rect 8660 -710 8860 -510
rect 8660 -1370 8860 -1170
rect 8660 -2030 8860 -1830
rect 8660 -2690 8860 -2490
rect 8660 -3350 8860 -3150
rect 6926 -4060 7126 -3860
rect 8660 -4010 8860 -3810
rect 8660 -4670 8860 -4470
rect 8660 -5330 8860 -5130
rect 8660 -5990 8860 -5790
rect 8660 -6650 8860 -6450
rect 8660 -7310 8860 -7110
rect 6936 -7630 7136 -7430
rect 8660 -7970 8860 -7770
rect 8660 -8630 8860 -8430
rect 8660 -9290 8860 -9090
rect 8660 -9950 8860 -9750
rect 7820 -10610 8020 -10410
rect 8660 -10610 8860 -10410
<< metal4 >>
rect 1330 1480 1470 1500
rect 1330 1380 1350 1480
rect 1450 1380 1470 1480
rect 1330 1360 1470 1380
rect 1350 -410 1450 1360
rect 8610 860 8910 930
rect 8610 660 8660 860
rect 8860 660 8910 860
rect 8610 150 8910 660
rect 8610 -50 8660 150
rect 8860 -50 8910 150
rect 8610 -510 8910 -50
rect 8610 -710 8660 -510
rect 8860 -710 8910 -510
rect 8610 -1170 8910 -710
rect 8610 -1370 8660 -1170
rect 8860 -1370 8910 -1170
rect 8610 -1830 8910 -1370
rect 8610 -2030 8660 -1830
rect 8860 -2030 8910 -1830
rect 8610 -2490 8910 -2030
rect 8610 -2690 8660 -2490
rect 8860 -2690 8910 -2490
rect 8610 -3150 8910 -2690
rect 8610 -3250 8660 -3150
rect 8170 -3350 8660 -3250
rect 8860 -3350 8910 -3150
rect 8170 -3550 8910 -3350
rect 8610 -3810 8910 -3550
rect 6906 -3860 7146 -3840
rect 6906 -4060 6926 -3860
rect 7126 -4060 7146 -3860
rect 6906 -4080 7146 -4060
rect 8610 -4010 8660 -3810
rect 8860 -4010 8910 -3810
rect 8610 -4470 8910 -4010
rect 8610 -4670 8660 -4470
rect 8860 -4670 8910 -4470
rect 8610 -5130 8910 -4670
rect 8610 -5330 8660 -5130
rect 8860 -5330 8910 -5130
rect 8610 -5790 8910 -5330
rect 8610 -5990 8660 -5790
rect 8860 -5990 8910 -5790
rect 8610 -6450 8910 -5990
rect 8610 -6650 8660 -6450
rect 8860 -6650 8910 -6450
rect 8610 -6790 8910 -6650
rect 8190 -7090 8910 -6790
rect 8610 -7110 8910 -7090
rect 8610 -7310 8660 -7110
rect 8860 -7310 8910 -7110
rect 6916 -7430 7156 -7410
rect 6916 -7630 6936 -7430
rect 7136 -7630 7156 -7430
rect 6916 -7650 7156 -7630
rect 8610 -7770 8910 -7310
rect 8610 -7970 8660 -7770
rect 8860 -7970 8910 -7770
rect 8610 -8430 8910 -7970
rect 8610 -8630 8660 -8430
rect 8860 -8630 8910 -8430
rect 8610 -9090 8910 -8630
rect 8610 -9290 8660 -9090
rect 8860 -9290 8910 -9090
rect 8610 -9750 8910 -9290
rect 8610 -9950 8660 -9750
rect 8860 -9950 8910 -9750
rect 8610 -10360 8910 -9950
rect 7770 -10410 8070 -10360
rect 7770 -10610 7820 -10410
rect 8020 -10610 8070 -10410
rect 7770 -10660 8070 -10610
rect 8190 -10410 8910 -10360
rect 8190 -10610 8660 -10410
rect 8860 -10610 8910 -10410
rect 8190 -10660 8910 -10610
use cbank  cbank_0
timestamp 1640901595
transform 1 0 -84 0 1 -1870
box -30 -1680 8150 1550
use cbank  cbank_2
timestamp 1640901595
transform 1 0 -84 0 1 -8980
box -30 -1680 8150 1550
use cbank  cbank_1
timestamp 1640901595
transform 1 0 -84 0 1 -5410
box -30 -1680 8150 1550
use ro_var_extend  ro_var_extend_0
timestamp 1640901061
transform 1 0 974 0 1 1350
box -250 -800 6290 1010
<< labels >>
rlabel locali 2246 -1650 2246 -1650 1 a0
rlabel locali 3234 -1660 3234 -1660 1 a1
rlabel locali 7346 -1650 7346 -1650 1 a5
rlabel locali 6144 -1650 6144 -1650 1 a4
rlabel locali 5182 -1650 5182 -1650 1 a3
rlabel locali 4202 -1670 4202 -1670 1 a2
<< end >>
