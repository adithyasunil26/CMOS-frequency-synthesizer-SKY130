magic
tech sky130A
timestamp 1640994530
<< locali >>
rect 225 3125 235 3145
rect 255 3125 275 3145
<< viali >>
rect 260 3635 280 3655
rect 235 3125 255 3145
rect 4865 645 4885 665
<< metal1 >>
rect 250 3655 290 3665
rect 175 3635 260 3655
rect 280 3635 290 3655
rect 175 2750 195 3635
rect 250 3625 290 3635
rect 225 3150 265 3155
rect 225 3120 230 3150
rect 260 3120 265 3150
rect 225 3115 265 3120
rect 165 2745 205 2750
rect 165 2715 170 2745
rect 200 2715 205 2745
rect 165 2710 205 2715
rect 7050 1205 7085 1215
rect 7005 1190 7085 1205
rect 7050 1180 7085 1190
rect 7055 1070 7090 1080
rect 7005 1055 7090 1070
rect 7055 1045 7090 1055
rect 4855 670 4895 675
rect 4855 640 4860 670
rect 4890 640 4895 670
rect 4855 635 4895 640
<< via1 >>
rect 230 3145 260 3150
rect 230 3125 235 3145
rect 235 3125 255 3145
rect 255 3125 260 3145
rect 230 3120 260 3125
rect 170 2715 200 2745
rect 4860 665 4890 670
rect 4860 645 4865 665
rect 4865 645 4885 665
rect 4885 645 4890 665
rect 4860 640 4890 645
<< metal2 >>
rect 220 3155 270 3160
rect 220 3115 225 3155
rect 265 3115 270 3155
rect 220 3110 270 3115
rect 160 2750 210 2755
rect 160 2710 165 2750
rect 205 2710 210 2750
rect 160 2705 210 2710
rect 730 2050 775 2055
rect 730 2015 735 2050
rect 770 2015 775 2050
rect 730 2010 775 2015
rect 5410 1240 5445 1275
rect 245 685 285 695
rect 245 665 315 685
rect 4850 670 4900 680
rect 245 655 285 665
rect 4850 640 4860 670
rect 4890 640 4900 670
rect 4850 630 4900 640
rect 5190 425 5240 435
rect 5190 395 5200 425
rect 5230 415 5240 425
rect 5230 400 5430 415
rect 5230 395 5240 400
rect 5190 385 5240 395
<< via2 >>
rect 225 3150 265 3155
rect 225 3120 230 3150
rect 230 3120 260 3150
rect 260 3120 265 3150
rect 225 3115 265 3120
rect 165 2745 205 2750
rect 165 2715 170 2745
rect 170 2715 200 2745
rect 200 2715 205 2745
rect 165 2710 205 2715
rect 735 2015 770 2050
rect 4860 640 4890 670
rect 5200 395 5230 425
<< metal3 >>
rect 215 3155 275 3165
rect 215 3115 225 3155
rect 265 3115 275 3155
rect 215 3105 275 3115
rect 160 2750 210 2755
rect 160 2710 165 2750
rect 205 2725 210 2750
rect 205 2710 4895 2725
rect 160 2705 4895 2710
rect 165 2695 4895 2705
rect 725 2050 780 2060
rect 725 2015 735 2050
rect 770 2015 780 2050
rect 725 2005 780 2015
rect 4855 680 4895 2695
rect 4850 670 4900 680
rect 4850 640 4860 670
rect 4890 640 4900 670
rect 4850 630 4900 640
rect 5190 430 5240 435
rect 5190 390 5195 430
rect 5235 390 5240 430
rect 5190 385 5240 390
<< via3 >>
rect 225 3115 265 3155
rect 735 2015 770 2050
rect 5195 425 5235 430
rect 5195 395 5200 425
rect 5200 395 5230 425
rect 5230 395 5235 425
rect 5195 390 5235 395
<< metal4 >>
rect 210 3155 280 3170
rect 210 3115 225 3155
rect 265 3115 280 3155
rect 210 3100 280 3115
rect 220 2475 265 3100
rect 220 2435 5230 2475
rect 745 2110 800 2150
rect 745 2060 775 2110
rect 725 2050 780 2060
rect 725 2015 735 2050
rect 770 2015 780 2050
rect 725 2005 780 2015
rect 5200 435 5230 2435
rect 5190 430 5240 435
rect 5190 390 5195 430
rect 5235 390 5240 430
rect 5190 385 5240 390
use pd  pd_0
timestamp 1640980777
transform 1 0 5535 0 1 855
box -215 -855 1685 810
use divbuf  divbuf_0
timestamp 1640994347
transform 1 0 460 0 1 3640
box -460 -1085 31200 495
use divider  divider_0
timestamp 1640980777
transform 1 0 490 0 1 235
box -490 -235 4690 2150
<< labels >>
rlabel metal2 5240 400 5305 415 1 div
rlabel space 220 3125 285 3145 1 div
rlabel metal4 220 2435 5230 2475 1 div
rlabel metal3 4855 635 4895 2175 1 bufin
rlabel metal1 175 2720 195 3655 1 bufin
<< end >>
